// scala

module MULADD_2 (
  input      [51:0]   src1,
  input      [33:0]   src2,
  output     [65:0]   result
);

endmodule