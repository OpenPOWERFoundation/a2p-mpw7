VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM128
  CLASS BLOCK ;
  FOREIGN RAM128 ;
  ORIGIN 0.000 0.000 ;
  SIZE 399.740 BY 394.400 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 397.740 180.240 399.740 180.840 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 397.740 213.560 399.740 214.160 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 397.740 246.200 399.740 246.800 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 397.740 278.840 399.740 279.440 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 397.740 312.160 399.740 312.760 ;
    END
  END A0[4]
  PIN A0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 397.740 344.800 399.740 345.400 ;
    END
  END A0[5]
  PIN A0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 397.740 377.440 399.740 378.040 ;
    END
  END A0[6]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 2.000 197.840 ;
    END
  END CLK
  PIN Di0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 0.000 6.350 2.000 ;
    END
  END Di0[0]
  PIN Di0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.730 0.000 131.010 2.000 ;
    END
  END Di0[10]
  PIN Di0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.150 0.000 143.430 2.000 ;
    END
  END Di0[11]
  PIN Di0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 0.000 155.850 2.000 ;
    END
  END Di0[12]
  PIN Di0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 0.000 168.730 2.000 ;
    END
  END Di0[13]
  PIN Di0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.870 0.000 181.150 2.000 ;
    END
  END Di0[14]
  PIN Di0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 2.000 ;
    END
  END Di0[15]
  PIN Di0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 0.000 205.990 2.000 ;
    END
  END Di0[16]
  PIN Di0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 0.000 218.410 2.000 ;
    END
  END Di0[17]
  PIN Di0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 0.000 230.830 2.000 ;
    END
  END Di0[18]
  PIN Di0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 0.000 243.250 2.000 ;
    END
  END Di0[19]
  PIN Di0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 2.000 ;
    END
  END Di0[1]
  PIN Di0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.850 0.000 256.130 2.000 ;
    END
  END Di0[20]
  PIN Di0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 0.000 268.550 2.000 ;
    END
  END Di0[21]
  PIN Di0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 0.000 280.970 2.000 ;
    END
  END Di0[22]
  PIN Di0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 2.000 ;
    END
  END Di0[23]
  PIN Di0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.530 0.000 305.810 2.000 ;
    END
  END Di0[24]
  PIN Di0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 0.000 318.230 2.000 ;
    END
  END Di0[25]
  PIN Di0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 0.000 331.110 2.000 ;
    END
  END Di0[26]
  PIN Di0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.250 0.000 343.530 2.000 ;
    END
  END Di0[27]
  PIN Di0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.670 0.000 355.950 2.000 ;
    END
  END Di0[28]
  PIN Di0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.090 0.000 368.370 2.000 ;
    END
  END Di0[29]
  PIN Di0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 2.000 ;
    END
  END Di0[2]
  PIN Di0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.510 0.000 380.790 2.000 ;
    END
  END Di0[30]
  PIN Di0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 2.000 ;
    END
  END Di0[31]
  PIN Di0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 2.000 ;
    END
  END Di0[3]
  PIN Di0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 2.000 ;
    END
  END Di0[4]
  PIN Di0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 2.000 ;
    END
  END Di0[5]
  PIN Di0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 2.000 ;
    END
  END Di0[6]
  PIN Di0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 2.000 ;
    END
  END Di0[7]
  PIN Di0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 2.000 ;
    END
  END Di0[8]
  PIN Di0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.310 0.000 118.590 2.000 ;
    END
  END Di0[9]
  PIN Do0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 392.400 6.350 394.400 ;
    END
  END Do0[0]
  PIN Do0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.730 392.400 131.010 394.400 ;
    END
  END Do0[10]
  PIN Do0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.150 392.400 143.430 394.400 ;
    END
  END Do0[11]
  PIN Do0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 392.400 155.850 394.400 ;
    END
  END Do0[12]
  PIN Do0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 392.400 168.730 394.400 ;
    END
  END Do0[13]
  PIN Do0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.870 392.400 181.150 394.400 ;
    END
  END Do0[14]
  PIN Do0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 392.400 193.570 394.400 ;
    END
  END Do0[15]
  PIN Do0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 392.400 205.990 394.400 ;
    END
  END Do0[16]
  PIN Do0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 392.400 218.410 394.400 ;
    END
  END Do0[17]
  PIN Do0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 392.400 230.830 394.400 ;
    END
  END Do0[18]
  PIN Do0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 392.400 243.250 394.400 ;
    END
  END Do0[19]
  PIN Do0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 392.400 18.770 394.400 ;
    END
  END Do0[1]
  PIN Do0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.850 392.400 256.130 394.400 ;
    END
  END Do0[20]
  PIN Do0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 392.400 268.550 394.400 ;
    END
  END Do0[21]
  PIN Do0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 392.400 280.970 394.400 ;
    END
  END Do0[22]
  PIN Do0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 392.400 293.390 394.400 ;
    END
  END Do0[23]
  PIN Do0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.530 392.400 305.810 394.400 ;
    END
  END Do0[24]
  PIN Do0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 392.400 318.230 394.400 ;
    END
  END Do0[25]
  PIN Do0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 392.400 331.110 394.400 ;
    END
  END Do0[26]
  PIN Do0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.250 392.400 343.530 394.400 ;
    END
  END Do0[27]
  PIN Do0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.670 392.400 355.950 394.400 ;
    END
  END Do0[28]
  PIN Do0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.090 392.400 368.370 394.400 ;
    END
  END Do0[29]
  PIN Do0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 392.400 31.190 394.400 ;
    END
  END Do0[2]
  PIN Do0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.510 392.400 380.790 394.400 ;
    END
  END Do0[30]
  PIN Do0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 392.400 393.210 394.400 ;
    END
  END Do0[31]
  PIN Do0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 392.400 43.610 394.400 ;
    END
  END Do0[3]
  PIN Do0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 392.400 56.030 394.400 ;
    END
  END Do0[4]
  PIN Do0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 392.400 68.450 394.400 ;
    END
  END Do0[5]
  PIN Do0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 392.400 80.870 394.400 ;
    END
  END Do0[6]
  PIN Do0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 392.400 93.750 394.400 ;
    END
  END Do0[7]
  PIN Do0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 392.400 106.170 394.400 ;
    END
  END Do0[8]
  PIN Do0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.310 392.400 118.590 394.400 ;
    END
  END Do0[9]
  PIN EN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 397.740 16.360 399.740 16.960 ;
    END
  END EN0
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 95.080 2.480 96.680 391.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 248.680 2.480 250.280 391.920 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 18.280 2.480 19.880 391.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.880 2.480 173.480 391.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.480 2.480 327.080 391.920 ;
    END
  END VPWR
  PIN WE0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 397.740 49.000 399.740 49.600 ;
    END
  END WE0[0]
  PIN WE0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 397.740 81.640 399.740 82.240 ;
    END
  END WE0[1]
  PIN WE0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 397.740 114.960 399.740 115.560 ;
    END
  END WE0[2]
  PIN WE0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 397.740 147.600 399.740 148.200 ;
    END
  END WE0[3]
  OBS
      LAYER li1 ;
        RECT 2.760 2.635 396.980 391.765 ;
      LAYER met1 ;
        RECT 2.760 0.720 399.670 394.360 ;
      LAYER met2 ;
        RECT 3.320 392.120 5.790 394.390 ;
        RECT 6.630 392.120 18.210 394.390 ;
        RECT 19.050 392.120 30.630 394.390 ;
        RECT 31.470 392.120 43.050 394.390 ;
        RECT 43.890 392.120 55.470 394.390 ;
        RECT 56.310 392.120 67.890 394.390 ;
        RECT 68.730 392.120 80.310 394.390 ;
        RECT 81.150 392.120 93.190 394.390 ;
        RECT 94.030 392.120 105.610 394.390 ;
        RECT 106.450 392.120 118.030 394.390 ;
        RECT 118.870 392.120 130.450 394.390 ;
        RECT 131.290 392.120 142.870 394.390 ;
        RECT 143.710 392.120 155.290 394.390 ;
        RECT 156.130 392.120 168.170 394.390 ;
        RECT 169.010 392.120 180.590 394.390 ;
        RECT 181.430 392.120 193.010 394.390 ;
        RECT 193.850 392.120 205.430 394.390 ;
        RECT 206.270 392.120 217.850 394.390 ;
        RECT 218.690 392.120 230.270 394.390 ;
        RECT 231.110 392.120 242.690 394.390 ;
        RECT 243.530 392.120 255.570 394.390 ;
        RECT 256.410 392.120 267.990 394.390 ;
        RECT 268.830 392.120 280.410 394.390 ;
        RECT 281.250 392.120 292.830 394.390 ;
        RECT 293.670 392.120 305.250 394.390 ;
        RECT 306.090 392.120 317.670 394.390 ;
        RECT 318.510 392.120 330.550 394.390 ;
        RECT 331.390 392.120 342.970 394.390 ;
        RECT 343.810 392.120 355.390 394.390 ;
        RECT 356.230 392.120 367.810 394.390 ;
        RECT 368.650 392.120 380.230 394.390 ;
        RECT 381.070 392.120 392.650 394.390 ;
        RECT 393.490 392.120 399.640 394.390 ;
        RECT 3.320 2.280 399.640 392.120 ;
        RECT 3.320 0.155 5.790 2.280 ;
        RECT 6.630 0.155 18.210 2.280 ;
        RECT 19.050 0.155 30.630 2.280 ;
        RECT 31.470 0.155 43.050 2.280 ;
        RECT 43.890 0.155 55.470 2.280 ;
        RECT 56.310 0.155 67.890 2.280 ;
        RECT 68.730 0.155 80.310 2.280 ;
        RECT 81.150 0.155 93.190 2.280 ;
        RECT 94.030 0.155 105.610 2.280 ;
        RECT 106.450 0.155 118.030 2.280 ;
        RECT 118.870 0.155 130.450 2.280 ;
        RECT 131.290 0.155 142.870 2.280 ;
        RECT 143.710 0.155 155.290 2.280 ;
        RECT 156.130 0.155 168.170 2.280 ;
        RECT 169.010 0.155 180.590 2.280 ;
        RECT 181.430 0.155 193.010 2.280 ;
        RECT 193.850 0.155 205.430 2.280 ;
        RECT 206.270 0.155 217.850 2.280 ;
        RECT 218.690 0.155 230.270 2.280 ;
        RECT 231.110 0.155 242.690 2.280 ;
        RECT 243.530 0.155 255.570 2.280 ;
        RECT 256.410 0.155 267.990 2.280 ;
        RECT 268.830 0.155 280.410 2.280 ;
        RECT 281.250 0.155 292.830 2.280 ;
        RECT 293.670 0.155 305.250 2.280 ;
        RECT 306.090 0.155 317.670 2.280 ;
        RECT 318.510 0.155 330.550 2.280 ;
        RECT 331.390 0.155 342.970 2.280 ;
        RECT 343.810 0.155 355.390 2.280 ;
        RECT 356.230 0.155 367.810 2.280 ;
        RECT 368.650 0.155 380.230 2.280 ;
        RECT 381.070 0.155 392.650 2.280 ;
        RECT 393.490 0.155 399.640 2.280 ;
      LAYER met3 ;
        RECT 2.000 378.440 397.835 394.225 ;
        RECT 2.000 377.040 397.340 378.440 ;
        RECT 2.000 345.800 397.835 377.040 ;
        RECT 2.000 344.400 397.340 345.800 ;
        RECT 2.000 313.160 397.835 344.400 ;
        RECT 2.000 311.760 397.340 313.160 ;
        RECT 2.000 279.840 397.835 311.760 ;
        RECT 2.000 278.440 397.340 279.840 ;
        RECT 2.000 247.200 397.835 278.440 ;
        RECT 2.000 245.800 397.340 247.200 ;
        RECT 2.000 214.560 397.835 245.800 ;
        RECT 2.000 213.160 397.340 214.560 ;
        RECT 2.000 198.240 397.835 213.160 ;
        RECT 2.400 196.840 397.835 198.240 ;
        RECT 2.000 181.240 397.835 196.840 ;
        RECT 2.000 179.840 397.340 181.240 ;
        RECT 2.000 148.600 397.835 179.840 ;
        RECT 2.000 147.200 397.340 148.600 ;
        RECT 2.000 115.960 397.835 147.200 ;
        RECT 2.000 114.560 397.340 115.960 ;
        RECT 2.000 82.640 397.835 114.560 ;
        RECT 2.000 81.240 397.340 82.640 ;
        RECT 2.000 50.000 397.835 81.240 ;
        RECT 2.000 48.600 397.340 50.000 ;
        RECT 2.000 17.360 397.835 48.600 ;
        RECT 2.000 15.960 397.340 17.360 ;
        RECT 2.000 0.175 397.835 15.960 ;
      LAYER met4 ;
        RECT 38.015 392.320 383.345 394.225 ;
        RECT 38.015 43.015 94.680 392.320 ;
        RECT 97.080 43.015 171.480 392.320 ;
        RECT 173.880 43.015 248.280 392.320 ;
        RECT 250.680 43.015 325.080 392.320 ;
        RECT 327.480 43.015 383.345 392.320 ;
  END
END RAM128
END LIBRARY

