// scala

module MULADD_1 (
  input      [32:0]   src1,
  input      [49:0]   src2,
  input      [49:0]   src3,
  output     [51:0]   result
);
endmodule