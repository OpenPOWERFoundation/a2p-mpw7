VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DFFRF_3R1W
  CLASS BLOCK ;
  FOREIGN DFFRF_3R1W ;
  ORIGIN 0.000 0.000 ;
  SIZE 495.880 BY 266.560 ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 2.000 133.240 ;
    END
  END CLK
  PIN DA[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 264.560 7.730 266.560 ;
    END
  END DA[0]
  PIN DA[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 264.560 58.330 266.560 ;
    END
  END DA[10]
  PIN DA[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 264.560 63.390 266.560 ;
    END
  END DA[11]
  PIN DA[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 264.560 68.450 266.560 ;
    END
  END DA[12]
  PIN DA[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 264.560 73.510 266.560 ;
    END
  END DA[13]
  PIN DA[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 264.560 78.570 266.560 ;
    END
  END DA[14]
  PIN DA[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 264.560 83.630 266.560 ;
    END
  END DA[15]
  PIN DA[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 264.560 88.690 266.560 ;
    END
  END DA[16]
  PIN DA[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 264.560 93.750 266.560 ;
    END
  END DA[17]
  PIN DA[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 264.560 98.810 266.560 ;
    END
  END DA[18]
  PIN DA[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 264.560 103.870 266.560 ;
    END
  END DA[19]
  PIN DA[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 264.560 12.790 266.560 ;
    END
  END DA[1]
  PIN DA[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 264.560 108.930 266.560 ;
    END
  END DA[20]
  PIN DA[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 264.560 113.990 266.560 ;
    END
  END DA[21]
  PIN DA[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 264.560 119.050 266.560 ;
    END
  END DA[22]
  PIN DA[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.830 264.560 124.110 266.560 ;
    END
  END DA[23]
  PIN DA[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 264.560 129.170 266.560 ;
    END
  END DA[24]
  PIN DA[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 264.560 134.230 266.560 ;
    END
  END DA[25]
  PIN DA[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 264.560 139.290 266.560 ;
    END
  END DA[26]
  PIN DA[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 264.560 144.350 266.560 ;
    END
  END DA[27]
  PIN DA[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 264.560 149.410 266.560 ;
    END
  END DA[28]
  PIN DA[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.190 264.560 154.470 266.560 ;
    END
  END DA[29]
  PIN DA[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 264.560 17.850 266.560 ;
    END
  END DA[2]
  PIN DA[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 264.560 159.530 266.560 ;
    END
  END DA[30]
  PIN DA[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 264.560 164.590 266.560 ;
    END
  END DA[31]
  PIN DA[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 264.560 22.910 266.560 ;
    END
  END DA[3]
  PIN DA[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 264.560 27.970 266.560 ;
    END
  END DA[4]
  PIN DA[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.750 264.560 33.030 266.560 ;
    END
  END DA[5]
  PIN DA[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 264.560 38.090 266.560 ;
    END
  END DA[6]
  PIN DA[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 264.560 43.150 266.560 ;
    END
  END DA[7]
  PIN DA[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 264.560 48.210 266.560 ;
    END
  END DA[8]
  PIN DA[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 264.560 53.270 266.560 ;
    END
  END DA[9]
  PIN DB[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 264.560 169.650 266.560 ;
    END
  END DB[0]
  PIN DB[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.970 264.560 220.250 266.560 ;
    END
  END DB[10]
  PIN DB[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 264.560 225.310 266.560 ;
    END
  END DB[11]
  PIN DB[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.090 264.560 230.370 266.560 ;
    END
  END DB[12]
  PIN DB[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 264.560 235.430 266.560 ;
    END
  END DB[13]
  PIN DB[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 264.560 240.490 266.560 ;
    END
  END DB[14]
  PIN DB[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.270 264.560 245.550 266.560 ;
    END
  END DB[15]
  PIN DB[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.330 264.560 250.610 266.560 ;
    END
  END DB[16]
  PIN DB[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 264.560 255.670 266.560 ;
    END
  END DB[17]
  PIN DB[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.450 264.560 260.730 266.560 ;
    END
  END DB[18]
  PIN DB[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.510 264.560 265.790 266.560 ;
    END
  END DB[19]
  PIN DB[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 264.560 174.710 266.560 ;
    END
  END DB[1]
  PIN DB[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 264.560 270.850 266.560 ;
    END
  END DB[20]
  PIN DB[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.630 264.560 275.910 266.560 ;
    END
  END DB[21]
  PIN DB[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 264.560 280.970 266.560 ;
    END
  END DB[22]
  PIN DB[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.750 264.560 286.030 266.560 ;
    END
  END DB[23]
  PIN DB[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.810 264.560 291.090 266.560 ;
    END
  END DB[24]
  PIN DB[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.870 264.560 296.150 266.560 ;
    END
  END DB[25]
  PIN DB[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.930 264.560 301.210 266.560 ;
    END
  END DB[26]
  PIN DB[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 264.560 306.270 266.560 ;
    END
  END DB[27]
  PIN DB[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.050 264.560 311.330 266.560 ;
    END
  END DB[28]
  PIN DB[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.110 264.560 316.390 266.560 ;
    END
  END DB[29]
  PIN DB[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 264.560 179.770 266.560 ;
    END
  END DB[2]
  PIN DB[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.170 264.560 321.450 266.560 ;
    END
  END DB[30]
  PIN DB[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.230 264.560 326.510 266.560 ;
    END
  END DB[31]
  PIN DB[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.550 264.560 184.830 266.560 ;
    END
  END DB[3]
  PIN DB[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 264.560 189.890 266.560 ;
    END
  END DB[4]
  PIN DB[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 264.560 194.950 266.560 ;
    END
  END DB[5]
  PIN DB[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 264.560 200.010 266.560 ;
    END
  END DB[6]
  PIN DB[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.790 264.560 205.070 266.560 ;
    END
  END DB[7]
  PIN DB[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 264.560 210.130 266.560 ;
    END
  END DB[8]
  PIN DB[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 264.560 215.190 266.560 ;
    END
  END DB[9]
  PIN DC[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.290 264.560 331.570 266.560 ;
    END
  END DC[0]
  PIN DC[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.890 264.560 382.170 266.560 ;
    END
  END DC[10]
  PIN DC[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.950 264.560 387.230 266.560 ;
    END
  END DC[11]
  PIN DC[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 264.560 392.290 266.560 ;
    END
  END DC[12]
  PIN DC[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.070 264.560 397.350 266.560 ;
    END
  END DC[13]
  PIN DC[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.130 264.560 402.410 266.560 ;
    END
  END DC[14]
  PIN DC[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.190 264.560 407.470 266.560 ;
    END
  END DC[15]
  PIN DC[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 264.560 412.530 266.560 ;
    END
  END DC[16]
  PIN DC[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.310 264.560 417.590 266.560 ;
    END
  END DC[17]
  PIN DC[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.370 264.560 422.650 266.560 ;
    END
  END DC[18]
  PIN DC[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.430 264.560 427.710 266.560 ;
    END
  END DC[19]
  PIN DC[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.350 264.560 336.630 266.560 ;
    END
  END DC[1]
  PIN DC[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.490 264.560 432.770 266.560 ;
    END
  END DC[20]
  PIN DC[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.550 264.560 437.830 266.560 ;
    END
  END DC[21]
  PIN DC[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.610 264.560 442.890 266.560 ;
    END
  END DC[22]
  PIN DC[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 264.560 447.950 266.560 ;
    END
  END DC[23]
  PIN DC[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.730 264.560 453.010 266.560 ;
    END
  END DC[24]
  PIN DC[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.790 264.560 458.070 266.560 ;
    END
  END DC[25]
  PIN DC[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.850 264.560 463.130 266.560 ;
    END
  END DC[26]
  PIN DC[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.910 264.560 468.190 266.560 ;
    END
  END DC[27]
  PIN DC[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.970 264.560 473.250 266.560 ;
    END
  END DC[28]
  PIN DC[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.030 264.560 478.310 266.560 ;
    END
  END DC[29]
  PIN DC[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 264.560 341.690 266.560 ;
    END
  END DC[2]
  PIN DC[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 264.560 483.370 266.560 ;
    END
  END DC[30]
  PIN DC[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.150 264.560 488.430 266.560 ;
    END
  END DC[31]
  PIN DC[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.470 264.560 346.750 266.560 ;
    END
  END DC[3]
  PIN DC[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.530 264.560 351.810 266.560 ;
    END
  END DC[4]
  PIN DC[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.590 264.560 356.870 266.560 ;
    END
  END DC[5]
  PIN DC[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.650 264.560 361.930 266.560 ;
    END
  END DC[6]
  PIN DC[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.710 264.560 366.990 266.560 ;
    END
  END DC[7]
  PIN DC[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.770 264.560 372.050 266.560 ;
    END
  END DC[8]
  PIN DC[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 264.560 377.110 266.560 ;
    END
  END DC[9]
  PIN DW[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 0.000 12.790 2.000 ;
    END
  END DW[0]
  PIN DW[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 2.000 ;
    END
  END DW[10]
  PIN DW[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 0.000 179.770 2.000 ;
    END
  END DW[11]
  PIN DW[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 0.000 194.950 2.000 ;
    END
  END DW[12]
  PIN DW[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 2.000 ;
    END
  END DW[13]
  PIN DW[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 0.000 225.310 2.000 ;
    END
  END DW[14]
  PIN DW[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 0.000 240.490 2.000 ;
    END
  END DW[15]
  PIN DW[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 0.000 255.670 2.000 ;
    END
  END DW[16]
  PIN DW[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 2.000 ;
    END
  END DW[17]
  PIN DW[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.750 0.000 286.030 2.000 ;
    END
  END DW[18]
  PIN DW[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.930 0.000 301.210 2.000 ;
    END
  END DW[19]
  PIN DW[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 2.000 ;
    END
  END DW[1]
  PIN DW[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.110 0.000 316.390 2.000 ;
    END
  END DW[20]
  PIN DW[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.290 0.000 331.570 2.000 ;
    END
  END DW[21]
  PIN DW[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.470 0.000 346.750 2.000 ;
    END
  END DW[22]
  PIN DW[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.650 0.000 361.930 2.000 ;
    END
  END DW[23]
  PIN DW[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 0.000 377.110 2.000 ;
    END
  END DW[24]
  PIN DW[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 0.000 392.290 2.000 ;
    END
  END DW[25]
  PIN DW[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.190 0.000 407.470 2.000 ;
    END
  END DW[26]
  PIN DW[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.370 0.000 422.650 2.000 ;
    END
  END DW[27]
  PIN DW[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.550 0.000 437.830 2.000 ;
    END
  END DW[28]
  PIN DW[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.730 0.000 453.010 2.000 ;
    END
  END DW[29]
  PIN DW[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 2.000 ;
    END
  END DW[2]
  PIN DW[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.910 0.000 468.190 2.000 ;
    END
  END DW[30]
  PIN DW[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 0.000 483.370 2.000 ;
    END
  END DW[31]
  PIN DW[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 2.000 ;
    END
  END DW[3]
  PIN DW[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 0.000 73.510 2.000 ;
    END
  END DW[4]
  PIN DW[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 2.000 ;
    END
  END DW[5]
  PIN DW[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 0.000 103.870 2.000 ;
    END
  END DW[6]
  PIN DW[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 2.000 ;
    END
  END DW[7]
  PIN DW[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 0.000 134.230 2.000 ;
    END
  END DW[8]
  PIN DW[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 0.000 149.410 2.000 ;
    END
  END DW[9]
  PIN RA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 493.880 8.880 495.880 9.480 ;
    END
  END RA[0]
  PIN RA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 493.880 26.560 495.880 27.160 ;
    END
  END RA[1]
  PIN RA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 493.880 44.240 495.880 44.840 ;
    END
  END RA[2]
  PIN RA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 493.880 61.920 495.880 62.520 ;
    END
  END RA[3]
  PIN RA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 493.880 79.600 495.880 80.200 ;
    END
  END RA[4]
  PIN RB[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 493.880 97.280 495.880 97.880 ;
    END
  END RB[0]
  PIN RB[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 493.880 114.960 495.880 115.560 ;
    END
  END RB[1]
  PIN RB[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 493.880 132.640 495.880 133.240 ;
    END
  END RB[2]
  PIN RB[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 493.880 150.320 495.880 150.920 ;
    END
  END RB[3]
  PIN RB[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 493.880 168.000 495.880 168.600 ;
    END
  END RB[4]
  PIN RC[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 493.880 185.680 495.880 186.280 ;
    END
  END RC[0]
  PIN RC[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 493.880 203.360 495.880 203.960 ;
    END
  END RC[1]
  PIN RC[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 493.880 221.040 495.880 221.640 ;
    END
  END RC[2]
  PIN RC[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 493.880 238.720 495.880 239.320 ;
    END
  END RC[3]
  PIN RC[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 493.880 256.400 495.880 257.000 ;
    END
  END RC[4]
  PIN RW[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 2.000 19.000 ;
    END
  END RW[0]
  PIN RW[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.480 2.000 57.080 ;
    END
  END RW[1]
  PIN RW[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 94.560 2.000 95.160 ;
    END
  END RW[2]
  PIN RW[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.800 2.000 209.400 ;
    END
  END RW[3]
  PIN RW[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.880 2.000 247.480 ;
    END
  END RW[4]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 95.080 2.480 96.680 264.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 248.680 2.480 250.280 264.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 402.280 2.480 403.880 264.080 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 18.280 2.480 19.880 264.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.880 2.480 173.480 264.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.480 2.480 327.080 264.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 479.080 2.480 480.680 264.080 ;
    END
  END VPWR
  PIN WE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.720 2.000 171.320 ;
    END
  END WE
  OBS
      LAYER li1 ;
        RECT 2.760 2.635 493.120 263.925 ;
      LAYER met1 ;
        RECT 0.990 0.040 494.430 266.520 ;
      LAYER met2 ;
        RECT 1.020 264.280 7.170 266.550 ;
        RECT 8.010 264.280 12.230 266.550 ;
        RECT 13.070 264.280 17.290 266.550 ;
        RECT 18.130 264.280 22.350 266.550 ;
        RECT 23.190 264.280 27.410 266.550 ;
        RECT 28.250 264.280 32.470 266.550 ;
        RECT 33.310 264.280 37.530 266.550 ;
        RECT 38.370 264.280 42.590 266.550 ;
        RECT 43.430 264.280 47.650 266.550 ;
        RECT 48.490 264.280 52.710 266.550 ;
        RECT 53.550 264.280 57.770 266.550 ;
        RECT 58.610 264.280 62.830 266.550 ;
        RECT 63.670 264.280 67.890 266.550 ;
        RECT 68.730 264.280 72.950 266.550 ;
        RECT 73.790 264.280 78.010 266.550 ;
        RECT 78.850 264.280 83.070 266.550 ;
        RECT 83.910 264.280 88.130 266.550 ;
        RECT 88.970 264.280 93.190 266.550 ;
        RECT 94.030 264.280 98.250 266.550 ;
        RECT 99.090 264.280 103.310 266.550 ;
        RECT 104.150 264.280 108.370 266.550 ;
        RECT 109.210 264.280 113.430 266.550 ;
        RECT 114.270 264.280 118.490 266.550 ;
        RECT 119.330 264.280 123.550 266.550 ;
        RECT 124.390 264.280 128.610 266.550 ;
        RECT 129.450 264.280 133.670 266.550 ;
        RECT 134.510 264.280 138.730 266.550 ;
        RECT 139.570 264.280 143.790 266.550 ;
        RECT 144.630 264.280 148.850 266.550 ;
        RECT 149.690 264.280 153.910 266.550 ;
        RECT 154.750 264.280 158.970 266.550 ;
        RECT 159.810 264.280 164.030 266.550 ;
        RECT 164.870 264.280 169.090 266.550 ;
        RECT 169.930 264.280 174.150 266.550 ;
        RECT 174.990 264.280 179.210 266.550 ;
        RECT 180.050 264.280 184.270 266.550 ;
        RECT 185.110 264.280 189.330 266.550 ;
        RECT 190.170 264.280 194.390 266.550 ;
        RECT 195.230 264.280 199.450 266.550 ;
        RECT 200.290 264.280 204.510 266.550 ;
        RECT 205.350 264.280 209.570 266.550 ;
        RECT 210.410 264.280 214.630 266.550 ;
        RECT 215.470 264.280 219.690 266.550 ;
        RECT 220.530 264.280 224.750 266.550 ;
        RECT 225.590 264.280 229.810 266.550 ;
        RECT 230.650 264.280 234.870 266.550 ;
        RECT 235.710 264.280 239.930 266.550 ;
        RECT 240.770 264.280 244.990 266.550 ;
        RECT 245.830 264.280 250.050 266.550 ;
        RECT 250.890 264.280 255.110 266.550 ;
        RECT 255.950 264.280 260.170 266.550 ;
        RECT 261.010 264.280 265.230 266.550 ;
        RECT 266.070 264.280 270.290 266.550 ;
        RECT 271.130 264.280 275.350 266.550 ;
        RECT 276.190 264.280 280.410 266.550 ;
        RECT 281.250 264.280 285.470 266.550 ;
        RECT 286.310 264.280 290.530 266.550 ;
        RECT 291.370 264.280 295.590 266.550 ;
        RECT 296.430 264.280 300.650 266.550 ;
        RECT 301.490 264.280 305.710 266.550 ;
        RECT 306.550 264.280 310.770 266.550 ;
        RECT 311.610 264.280 315.830 266.550 ;
        RECT 316.670 264.280 320.890 266.550 ;
        RECT 321.730 264.280 325.950 266.550 ;
        RECT 326.790 264.280 331.010 266.550 ;
        RECT 331.850 264.280 336.070 266.550 ;
        RECT 336.910 264.280 341.130 266.550 ;
        RECT 341.970 264.280 346.190 266.550 ;
        RECT 347.030 264.280 351.250 266.550 ;
        RECT 352.090 264.280 356.310 266.550 ;
        RECT 357.150 264.280 361.370 266.550 ;
        RECT 362.210 264.280 366.430 266.550 ;
        RECT 367.270 264.280 371.490 266.550 ;
        RECT 372.330 264.280 376.550 266.550 ;
        RECT 377.390 264.280 381.610 266.550 ;
        RECT 382.450 264.280 386.670 266.550 ;
        RECT 387.510 264.280 391.730 266.550 ;
        RECT 392.570 264.280 396.790 266.550 ;
        RECT 397.630 264.280 401.850 266.550 ;
        RECT 402.690 264.280 406.910 266.550 ;
        RECT 407.750 264.280 411.970 266.550 ;
        RECT 412.810 264.280 417.030 266.550 ;
        RECT 417.870 264.280 422.090 266.550 ;
        RECT 422.930 264.280 427.150 266.550 ;
        RECT 427.990 264.280 432.210 266.550 ;
        RECT 433.050 264.280 437.270 266.550 ;
        RECT 438.110 264.280 442.330 266.550 ;
        RECT 443.170 264.280 447.390 266.550 ;
        RECT 448.230 264.280 452.450 266.550 ;
        RECT 453.290 264.280 457.510 266.550 ;
        RECT 458.350 264.280 462.570 266.550 ;
        RECT 463.410 264.280 467.630 266.550 ;
        RECT 468.470 264.280 472.690 266.550 ;
        RECT 473.530 264.280 477.750 266.550 ;
        RECT 478.590 264.280 482.810 266.550 ;
        RECT 483.650 264.280 487.870 266.550 ;
        RECT 488.710 264.280 494.400 266.550 ;
        RECT 1.020 2.280 494.400 264.280 ;
        RECT 1.020 0.010 12.230 2.280 ;
        RECT 13.070 0.010 27.410 2.280 ;
        RECT 28.250 0.010 42.590 2.280 ;
        RECT 43.430 0.010 57.770 2.280 ;
        RECT 58.610 0.010 72.950 2.280 ;
        RECT 73.790 0.010 88.130 2.280 ;
        RECT 88.970 0.010 103.310 2.280 ;
        RECT 104.150 0.010 118.490 2.280 ;
        RECT 119.330 0.010 133.670 2.280 ;
        RECT 134.510 0.010 148.850 2.280 ;
        RECT 149.690 0.010 164.030 2.280 ;
        RECT 164.870 0.010 179.210 2.280 ;
        RECT 180.050 0.010 194.390 2.280 ;
        RECT 195.230 0.010 209.570 2.280 ;
        RECT 210.410 0.010 224.750 2.280 ;
        RECT 225.590 0.010 239.930 2.280 ;
        RECT 240.770 0.010 255.110 2.280 ;
        RECT 255.950 0.010 270.290 2.280 ;
        RECT 271.130 0.010 285.470 2.280 ;
        RECT 286.310 0.010 300.650 2.280 ;
        RECT 301.490 0.010 315.830 2.280 ;
        RECT 316.670 0.010 331.010 2.280 ;
        RECT 331.850 0.010 346.190 2.280 ;
        RECT 347.030 0.010 361.370 2.280 ;
        RECT 362.210 0.010 376.550 2.280 ;
        RECT 377.390 0.010 391.730 2.280 ;
        RECT 392.570 0.010 406.910 2.280 ;
        RECT 407.750 0.010 422.090 2.280 ;
        RECT 422.930 0.010 437.270 2.280 ;
        RECT 438.110 0.010 452.450 2.280 ;
        RECT 453.290 0.010 467.630 2.280 ;
        RECT 468.470 0.010 482.810 2.280 ;
        RECT 483.650 0.010 494.400 2.280 ;
      LAYER met3 ;
        RECT 2.000 257.400 493.880 266.385 ;
        RECT 2.000 256.000 493.480 257.400 ;
        RECT 2.000 247.880 493.880 256.000 ;
        RECT 2.400 246.480 493.880 247.880 ;
        RECT 2.000 239.720 493.880 246.480 ;
        RECT 2.000 238.320 493.480 239.720 ;
        RECT 2.000 222.040 493.880 238.320 ;
        RECT 2.000 220.640 493.480 222.040 ;
        RECT 2.000 209.800 493.880 220.640 ;
        RECT 2.400 208.400 493.880 209.800 ;
        RECT 2.000 204.360 493.880 208.400 ;
        RECT 2.000 202.960 493.480 204.360 ;
        RECT 2.000 186.680 493.880 202.960 ;
        RECT 2.000 185.280 493.480 186.680 ;
        RECT 2.000 171.720 493.880 185.280 ;
        RECT 2.400 170.320 493.880 171.720 ;
        RECT 2.000 169.000 493.880 170.320 ;
        RECT 2.000 167.600 493.480 169.000 ;
        RECT 2.000 151.320 493.880 167.600 ;
        RECT 2.000 149.920 493.480 151.320 ;
        RECT 2.000 133.640 493.880 149.920 ;
        RECT 2.400 132.240 493.480 133.640 ;
        RECT 2.000 115.960 493.880 132.240 ;
        RECT 2.000 114.560 493.480 115.960 ;
        RECT 2.000 98.280 493.880 114.560 ;
        RECT 2.000 96.880 493.480 98.280 ;
        RECT 2.000 95.560 493.880 96.880 ;
        RECT 2.400 94.160 493.880 95.560 ;
        RECT 2.000 80.600 493.880 94.160 ;
        RECT 2.000 79.200 493.480 80.600 ;
        RECT 2.000 62.920 493.880 79.200 ;
        RECT 2.000 61.520 493.480 62.920 ;
        RECT 2.000 57.480 493.880 61.520 ;
        RECT 2.400 56.080 493.880 57.480 ;
        RECT 2.000 45.240 493.880 56.080 ;
        RECT 2.000 43.840 493.480 45.240 ;
        RECT 2.000 27.560 493.880 43.840 ;
        RECT 2.000 26.160 493.480 27.560 ;
        RECT 2.000 19.400 493.880 26.160 ;
        RECT 2.400 18.000 493.880 19.400 ;
        RECT 2.000 9.880 493.880 18.000 ;
        RECT 2.000 8.480 493.480 9.880 ;
        RECT 2.000 0.175 493.880 8.480 ;
      LAYER met4 ;
        RECT 3.055 13.095 17.880 256.865 ;
        RECT 20.280 13.095 94.680 256.865 ;
        RECT 97.080 13.095 171.480 256.865 ;
        RECT 173.880 13.095 248.280 256.865 ;
        RECT 250.680 13.095 325.080 256.865 ;
        RECT 327.480 13.095 401.880 256.865 ;
        RECT 404.280 13.095 478.680 256.865 ;
        RECT 481.080 13.095 481.785 256.865 ;
  END
END DFFRF_3R1W
END LIBRARY

