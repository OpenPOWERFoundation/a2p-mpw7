VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO GPR
  CLASS BLOCK ;
  FOREIGN GPR ;
  ORIGIN 0.000 0.000 ;
  SIZE 1000.000 BY 500.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 0.000 9.110 4.000 ;
    END
  END clk
  PIN rd_adr_0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.760 4.000 20.360 ;
    END
  END rd_adr_0[0]
  PIN rd_adr_0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END rd_adr_0[1]
  PIN rd_adr_0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 4.000 73.400 ;
    END
  END rd_adr_0[2]
  PIN rd_adr_0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END rd_adr_0[3]
  PIN rd_adr_0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END rd_adr_0[4]
  PIN rd_adr_1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END rd_adr_1[0]
  PIN rd_adr_1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.120 4.000 55.720 ;
    END
  END rd_adr_1[1]
  PIN rd_adr_1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END rd_adr_1[2]
  PIN rd_adr_1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.160 4.000 108.760 ;
    END
  END rd_adr_1[3]
  PIN rd_adr_1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 4.000 135.280 ;
    END
  END rd_adr_1[4]
  PIN rd_adr_2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END rd_adr_2[0]
  PIN rd_adr_2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END rd_adr_2[1]
  PIN rd_adr_2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 90.480 4.000 91.080 ;
    END
  END rd_adr_2[2]
  PIN rd_adr_2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END rd_adr_2[3]
  PIN rd_adr_2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 143.520 4.000 144.120 ;
    END
  END rd_adr_2[4]
  PIN rd_dat_0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END rd_dat_0[0]
  PIN rd_dat_0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.670 0.000 332.950 4.000 ;
    END
  END rd_dat_0[10]
  PIN rd_dat_0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.030 0.000 363.310 4.000 ;
    END
  END rd_dat_0[11]
  PIN rd_dat_0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.390 0.000 393.670 4.000 ;
    END
  END rd_dat_0[12]
  PIN rd_dat_0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.750 0.000 424.030 4.000 ;
    END
  END rd_dat_0[13]
  PIN rd_dat_0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 4.000 ;
    END
  END rd_dat_0[14]
  PIN rd_dat_0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.470 0.000 484.750 4.000 ;
    END
  END rd_dat_0[15]
  PIN rd_dat_0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.830 0.000 515.110 4.000 ;
    END
  END rd_dat_0[16]
  PIN rd_dat_0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.190 0.000 545.470 4.000 ;
    END
  END rd_dat_0[17]
  PIN rd_dat_0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.550 0.000 575.830 4.000 ;
    END
  END rd_dat_0[18]
  PIN rd_dat_0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.910 0.000 606.190 4.000 ;
    END
  END rd_dat_0[19]
  PIN rd_dat_0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 4.000 ;
    END
  END rd_dat_0[1]
  PIN rd_dat_0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.270 0.000 636.550 4.000 ;
    END
  END rd_dat_0[20]
  PIN rd_dat_0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.630 0.000 666.910 4.000 ;
    END
  END rd_dat_0[21]
  PIN rd_dat_0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.990 0.000 697.270 4.000 ;
    END
  END rd_dat_0[22]
  PIN rd_dat_0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.350 0.000 727.630 4.000 ;
    END
  END rd_dat_0[23]
  PIN rd_dat_0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.710 0.000 757.990 4.000 ;
    END
  END rd_dat_0[24]
  PIN rd_dat_0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.070 0.000 788.350 4.000 ;
    END
  END rd_dat_0[25]
  PIN rd_dat_0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.430 0.000 818.710 4.000 ;
    END
  END rd_dat_0[26]
  PIN rd_dat_0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 848.790 0.000 849.070 4.000 ;
    END
  END rd_dat_0[27]
  PIN rd_dat_0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.150 0.000 879.430 4.000 ;
    END
  END rd_dat_0[28]
  PIN rd_dat_0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.510 0.000 909.790 4.000 ;
    END
  END rd_dat_0[29]
  PIN rd_dat_0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 4.000 ;
    END
  END rd_dat_0[2]
  PIN rd_dat_0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 939.870 0.000 940.150 4.000 ;
    END
  END rd_dat_0[30]
  PIN rd_dat_0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 970.230 0.000 970.510 4.000 ;
    END
  END rd_dat_0[31]
  PIN rd_dat_0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 0.000 120.430 4.000 ;
    END
  END rd_dat_0[3]
  PIN rd_dat_0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 0.000 150.790 4.000 ;
    END
  END rd_dat_0[4]
  PIN rd_dat_0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.870 0.000 181.150 4.000 ;
    END
  END rd_dat_0[5]
  PIN rd_dat_0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 0.000 211.510 4.000 ;
    END
  END rd_dat_0[6]
  PIN rd_dat_0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END rd_dat_0[7]
  PIN rd_dat_0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.950 0.000 272.230 4.000 ;
    END
  END rd_dat_0[8]
  PIN rd_dat_0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 0.000 302.590 4.000 ;
    END
  END rd_dat_0[9]
  PIN rd_dat_1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 4.000 ;
    END
  END rd_dat_1[0]
  PIN rd_dat_1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 0.000 343.070 4.000 ;
    END
  END rd_dat_1[10]
  PIN rd_dat_1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.150 0.000 373.430 4.000 ;
    END
  END rd_dat_1[11]
  PIN rd_dat_1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.510 0.000 403.790 4.000 ;
    END
  END rd_dat_1[12]
  PIN rd_dat_1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.870 0.000 434.150 4.000 ;
    END
  END rd_dat_1[13]
  PIN rd_dat_1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.230 0.000 464.510 4.000 ;
    END
  END rd_dat_1[14]
  PIN rd_dat_1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.590 0.000 494.870 4.000 ;
    END
  END rd_dat_1[15]
  PIN rd_dat_1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 0.000 525.230 4.000 ;
    END
  END rd_dat_1[16]
  PIN rd_dat_1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.310 0.000 555.590 4.000 ;
    END
  END rd_dat_1[17]
  PIN rd_dat_1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.670 0.000 585.950 4.000 ;
    END
  END rd_dat_1[18]
  PIN rd_dat_1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.030 0.000 616.310 4.000 ;
    END
  END rd_dat_1[19]
  PIN rd_dat_1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 4.000 ;
    END
  END rd_dat_1[1]
  PIN rd_dat_1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.390 0.000 646.670 4.000 ;
    END
  END rd_dat_1[20]
  PIN rd_dat_1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.750 0.000 677.030 4.000 ;
    END
  END rd_dat_1[21]
  PIN rd_dat_1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.110 0.000 707.390 4.000 ;
    END
  END rd_dat_1[22]
  PIN rd_dat_1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.470 0.000 737.750 4.000 ;
    END
  END rd_dat_1[23]
  PIN rd_dat_1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.830 0.000 768.110 4.000 ;
    END
  END rd_dat_1[24]
  PIN rd_dat_1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.190 0.000 798.470 4.000 ;
    END
  END rd_dat_1[25]
  PIN rd_dat_1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.550 0.000 828.830 4.000 ;
    END
  END rd_dat_1[26]
  PIN rd_dat_1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 858.910 0.000 859.190 4.000 ;
    END
  END rd_dat_1[27]
  PIN rd_dat_1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.270 0.000 889.550 4.000 ;
    END
  END rd_dat_1[28]
  PIN rd_dat_1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 919.630 0.000 919.910 4.000 ;
    END
  END rd_dat_1[29]
  PIN rd_dat_1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END rd_dat_1[2]
  PIN rd_dat_1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.990 0.000 950.270 4.000 ;
    END
  END rd_dat_1[30]
  PIN rd_dat_1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 980.350 0.000 980.630 4.000 ;
    END
  END rd_dat_1[31]
  PIN rd_dat_1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 0.000 130.550 4.000 ;
    END
  END rd_dat_1[3]
  PIN rd_dat_1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.630 0.000 160.910 4.000 ;
    END
  END rd_dat_1[4]
  PIN rd_dat_1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 0.000 191.270 4.000 ;
    END
  END rd_dat_1[5]
  PIN rd_dat_1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.350 0.000 221.630 4.000 ;
    END
  END rd_dat_1[6]
  PIN rd_dat_1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.710 0.000 251.990 4.000 ;
    END
  END rd_dat_1[7]
  PIN rd_dat_1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.070 0.000 282.350 4.000 ;
    END
  END rd_dat_1[8]
  PIN rd_dat_1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 0.000 312.710 4.000 ;
    END
  END rd_dat_1[9]
  PIN rd_dat_2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 0.000 49.590 4.000 ;
    END
  END rd_dat_2[0]
  PIN rd_dat_2[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.910 0.000 353.190 4.000 ;
    END
  END rd_dat_2[10]
  PIN rd_dat_2[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 0.000 383.550 4.000 ;
    END
  END rd_dat_2[11]
  PIN rd_dat_2[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.630 0.000 413.910 4.000 ;
    END
  END rd_dat_2[12]
  PIN rd_dat_2[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.990 0.000 444.270 4.000 ;
    END
  END rd_dat_2[13]
  PIN rd_dat_2[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.350 0.000 474.630 4.000 ;
    END
  END rd_dat_2[14]
  PIN rd_dat_2[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.710 0.000 504.990 4.000 ;
    END
  END rd_dat_2[15]
  PIN rd_dat_2[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.070 0.000 535.350 4.000 ;
    END
  END rd_dat_2[16]
  PIN rd_dat_2[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.430 0.000 565.710 4.000 ;
    END
  END rd_dat_2[17]
  PIN rd_dat_2[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 0.000 596.070 4.000 ;
    END
  END rd_dat_2[18]
  PIN rd_dat_2[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.150 0.000 626.430 4.000 ;
    END
  END rd_dat_2[19]
  PIN rd_dat_2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 0.000 79.950 4.000 ;
    END
  END rd_dat_2[1]
  PIN rd_dat_2[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.510 0.000 656.790 4.000 ;
    END
  END rd_dat_2[20]
  PIN rd_dat_2[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.870 0.000 687.150 4.000 ;
    END
  END rd_dat_2[21]
  PIN rd_dat_2[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.230 0.000 717.510 4.000 ;
    END
  END rd_dat_2[22]
  PIN rd_dat_2[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.590 0.000 747.870 4.000 ;
    END
  END rd_dat_2[23]
  PIN rd_dat_2[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.950 0.000 778.230 4.000 ;
    END
  END rd_dat_2[24]
  PIN rd_dat_2[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.310 0.000 808.590 4.000 ;
    END
  END rd_dat_2[25]
  PIN rd_dat_2[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 838.670 0.000 838.950 4.000 ;
    END
  END rd_dat_2[26]
  PIN rd_dat_2[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.030 0.000 869.310 4.000 ;
    END
  END rd_dat_2[27]
  PIN rd_dat_2[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.390 0.000 899.670 4.000 ;
    END
  END rd_dat_2[28]
  PIN rd_dat_2[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 929.750 0.000 930.030 4.000 ;
    END
  END rd_dat_2[29]
  PIN rd_dat_2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 0.000 110.310 4.000 ;
    END
  END rd_dat_2[2]
  PIN rd_dat_2[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 960.110 0.000 960.390 4.000 ;
    END
  END rd_dat_2[30]
  PIN rd_dat_2[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 990.470 0.000 990.750 4.000 ;
    END
  END rd_dat_2[31]
  PIN rd_dat_2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 0.000 140.670 4.000 ;
    END
  END rd_dat_2[3]
  PIN rd_dat_2[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END rd_dat_2[4]
  PIN rd_dat_2[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.110 0.000 201.390 4.000 ;
    END
  END rd_dat_2[5]
  PIN rd_dat_2[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.470 0.000 231.750 4.000 ;
    END
  END rd_dat_2[6]
  PIN rd_dat_2[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 0.000 262.110 4.000 ;
    END
  END rd_dat_2[7]
  PIN rd_dat_2[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 0.000 292.470 4.000 ;
    END
  END rd_dat_2[8]
  PIN rd_dat_2[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 0.000 322.830 4.000 ;
    END
  END rd_dat_2[9]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 0.000 19.230 4.000 ;
    END
  END reset
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 487.120 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 487.120 ;
    END
  END vssd1
  PIN wr_adr_0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END wr_adr_0[0]
  PIN wr_adr_0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.200 4.000 161.800 ;
    END
  END wr_adr_0[1]
  PIN wr_adr_0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END wr_adr_0[2]
  PIN wr_adr_0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.880 4.000 179.480 ;
    END
  END wr_adr_0[3]
  PIN wr_adr_0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 4.000 188.320 ;
    END
  END wr_adr_0[4]
  PIN wr_dat_0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.560 4.000 197.160 ;
    END
  END wr_dat_0[0]
  PIN wr_dat_0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.960 4.000 285.560 ;
    END
  END wr_dat_0[10]
  PIN wr_dat_0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.800 4.000 294.400 ;
    END
  END wr_dat_0[11]
  PIN wr_dat_0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 302.640 4.000 303.240 ;
    END
  END wr_dat_0[12]
  PIN wr_dat_0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 311.480 4.000 312.080 ;
    END
  END wr_dat_0[13]
  PIN wr_dat_0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 320.320 4.000 320.920 ;
    END
  END wr_dat_0[14]
  PIN wr_dat_0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.160 4.000 329.760 ;
    END
  END wr_dat_0[15]
  PIN wr_dat_0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.000 4.000 338.600 ;
    END
  END wr_dat_0[16]
  PIN wr_dat_0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END wr_dat_0[17]
  PIN wr_dat_0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.680 4.000 356.280 ;
    END
  END wr_dat_0[18]
  PIN wr_dat_0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 364.520 4.000 365.120 ;
    END
  END wr_dat_0[19]
  PIN wr_dat_0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 4.000 206.000 ;
    END
  END wr_dat_0[1]
  PIN wr_dat_0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 373.360 4.000 373.960 ;
    END
  END wr_dat_0[20]
  PIN wr_dat_0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.200 4.000 382.800 ;
    END
  END wr_dat_0[21]
  PIN wr_dat_0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END wr_dat_0[22]
  PIN wr_dat_0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 399.880 4.000 400.480 ;
    END
  END wr_dat_0[23]
  PIN wr_dat_0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.720 4.000 409.320 ;
    END
  END wr_dat_0[24]
  PIN wr_dat_0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 417.560 4.000 418.160 ;
    END
  END wr_dat_0[25]
  PIN wr_dat_0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 426.400 4.000 427.000 ;
    END
  END wr_dat_0[26]
  PIN wr_dat_0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END wr_dat_0[27]
  PIN wr_dat_0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.080 4.000 444.680 ;
    END
  END wr_dat_0[28]
  PIN wr_dat_0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.920 4.000 453.520 ;
    END
  END wr_dat_0[29]
  PIN wr_dat_0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END wr_dat_0[2]
  PIN wr_dat_0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 461.760 4.000 462.360 ;
    END
  END wr_dat_0[30]
  PIN wr_dat_0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 470.600 4.000 471.200 ;
    END
  END wr_dat_0[31]
  PIN wr_dat_0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END wr_dat_0[3]
  PIN wr_dat_0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.920 4.000 232.520 ;
    END
  END wr_dat_0[4]
  PIN wr_dat_0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 4.000 241.360 ;
    END
  END wr_dat_0[5]
  PIN wr_dat_0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 249.600 4.000 250.200 ;
    END
  END wr_dat_0[6]
  PIN wr_dat_0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END wr_dat_0[7]
  PIN wr_dat_0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.280 4.000 267.880 ;
    END
  END wr_dat_0[8]
  PIN wr_dat_0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.120 4.000 276.720 ;
    END
  END wr_dat_0[9]
  PIN wr_en_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 479.440 4.000 480.040 ;
    END
  END wr_en_0
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 994.060 486.965 ;
      LAYER met1 ;
        RECT 5.520 0.040 994.060 487.120 ;
      LAYER met2 ;
        RECT 7.460 4.280 990.680 487.065 ;
        RECT 7.460 0.010 8.550 4.280 ;
        RECT 9.390 0.010 18.670 4.280 ;
        RECT 19.510 0.010 28.790 4.280 ;
        RECT 29.630 0.010 38.910 4.280 ;
        RECT 39.750 0.010 49.030 4.280 ;
        RECT 49.870 0.010 59.150 4.280 ;
        RECT 59.990 0.010 69.270 4.280 ;
        RECT 70.110 0.010 79.390 4.280 ;
        RECT 80.230 0.010 89.510 4.280 ;
        RECT 90.350 0.010 99.630 4.280 ;
        RECT 100.470 0.010 109.750 4.280 ;
        RECT 110.590 0.010 119.870 4.280 ;
        RECT 120.710 0.010 129.990 4.280 ;
        RECT 130.830 0.010 140.110 4.280 ;
        RECT 140.950 0.010 150.230 4.280 ;
        RECT 151.070 0.010 160.350 4.280 ;
        RECT 161.190 0.010 170.470 4.280 ;
        RECT 171.310 0.010 180.590 4.280 ;
        RECT 181.430 0.010 190.710 4.280 ;
        RECT 191.550 0.010 200.830 4.280 ;
        RECT 201.670 0.010 210.950 4.280 ;
        RECT 211.790 0.010 221.070 4.280 ;
        RECT 221.910 0.010 231.190 4.280 ;
        RECT 232.030 0.010 241.310 4.280 ;
        RECT 242.150 0.010 251.430 4.280 ;
        RECT 252.270 0.010 261.550 4.280 ;
        RECT 262.390 0.010 271.670 4.280 ;
        RECT 272.510 0.010 281.790 4.280 ;
        RECT 282.630 0.010 291.910 4.280 ;
        RECT 292.750 0.010 302.030 4.280 ;
        RECT 302.870 0.010 312.150 4.280 ;
        RECT 312.990 0.010 322.270 4.280 ;
        RECT 323.110 0.010 332.390 4.280 ;
        RECT 333.230 0.010 342.510 4.280 ;
        RECT 343.350 0.010 352.630 4.280 ;
        RECT 353.470 0.010 362.750 4.280 ;
        RECT 363.590 0.010 372.870 4.280 ;
        RECT 373.710 0.010 382.990 4.280 ;
        RECT 383.830 0.010 393.110 4.280 ;
        RECT 393.950 0.010 403.230 4.280 ;
        RECT 404.070 0.010 413.350 4.280 ;
        RECT 414.190 0.010 423.470 4.280 ;
        RECT 424.310 0.010 433.590 4.280 ;
        RECT 434.430 0.010 443.710 4.280 ;
        RECT 444.550 0.010 453.830 4.280 ;
        RECT 454.670 0.010 463.950 4.280 ;
        RECT 464.790 0.010 474.070 4.280 ;
        RECT 474.910 0.010 484.190 4.280 ;
        RECT 485.030 0.010 494.310 4.280 ;
        RECT 495.150 0.010 504.430 4.280 ;
        RECT 505.270 0.010 514.550 4.280 ;
        RECT 515.390 0.010 524.670 4.280 ;
        RECT 525.510 0.010 534.790 4.280 ;
        RECT 535.630 0.010 544.910 4.280 ;
        RECT 545.750 0.010 555.030 4.280 ;
        RECT 555.870 0.010 565.150 4.280 ;
        RECT 565.990 0.010 575.270 4.280 ;
        RECT 576.110 0.010 585.390 4.280 ;
        RECT 586.230 0.010 595.510 4.280 ;
        RECT 596.350 0.010 605.630 4.280 ;
        RECT 606.470 0.010 615.750 4.280 ;
        RECT 616.590 0.010 625.870 4.280 ;
        RECT 626.710 0.010 635.990 4.280 ;
        RECT 636.830 0.010 646.110 4.280 ;
        RECT 646.950 0.010 656.230 4.280 ;
        RECT 657.070 0.010 666.350 4.280 ;
        RECT 667.190 0.010 676.470 4.280 ;
        RECT 677.310 0.010 686.590 4.280 ;
        RECT 687.430 0.010 696.710 4.280 ;
        RECT 697.550 0.010 706.830 4.280 ;
        RECT 707.670 0.010 716.950 4.280 ;
        RECT 717.790 0.010 727.070 4.280 ;
        RECT 727.910 0.010 737.190 4.280 ;
        RECT 738.030 0.010 747.310 4.280 ;
        RECT 748.150 0.010 757.430 4.280 ;
        RECT 758.270 0.010 767.550 4.280 ;
        RECT 768.390 0.010 777.670 4.280 ;
        RECT 778.510 0.010 787.790 4.280 ;
        RECT 788.630 0.010 797.910 4.280 ;
        RECT 798.750 0.010 808.030 4.280 ;
        RECT 808.870 0.010 818.150 4.280 ;
        RECT 818.990 0.010 828.270 4.280 ;
        RECT 829.110 0.010 838.390 4.280 ;
        RECT 839.230 0.010 848.510 4.280 ;
        RECT 849.350 0.010 858.630 4.280 ;
        RECT 859.470 0.010 868.750 4.280 ;
        RECT 869.590 0.010 878.870 4.280 ;
        RECT 879.710 0.010 888.990 4.280 ;
        RECT 889.830 0.010 899.110 4.280 ;
        RECT 899.950 0.010 909.230 4.280 ;
        RECT 910.070 0.010 919.350 4.280 ;
        RECT 920.190 0.010 929.470 4.280 ;
        RECT 930.310 0.010 939.590 4.280 ;
        RECT 940.430 0.010 949.710 4.280 ;
        RECT 950.550 0.010 959.830 4.280 ;
        RECT 960.670 0.010 969.950 4.280 ;
        RECT 970.790 0.010 980.070 4.280 ;
        RECT 980.910 0.010 990.190 4.280 ;
      LAYER met3 ;
        RECT 3.070 480.440 966.395 487.045 ;
        RECT 4.400 479.040 966.395 480.440 ;
        RECT 3.070 471.600 966.395 479.040 ;
        RECT 4.400 470.200 966.395 471.600 ;
        RECT 3.070 462.760 966.395 470.200 ;
        RECT 4.400 461.360 966.395 462.760 ;
        RECT 3.070 453.920 966.395 461.360 ;
        RECT 4.400 452.520 966.395 453.920 ;
        RECT 3.070 445.080 966.395 452.520 ;
        RECT 4.400 443.680 966.395 445.080 ;
        RECT 3.070 436.240 966.395 443.680 ;
        RECT 4.400 434.840 966.395 436.240 ;
        RECT 3.070 427.400 966.395 434.840 ;
        RECT 4.400 426.000 966.395 427.400 ;
        RECT 3.070 418.560 966.395 426.000 ;
        RECT 4.400 417.160 966.395 418.560 ;
        RECT 3.070 409.720 966.395 417.160 ;
        RECT 4.400 408.320 966.395 409.720 ;
        RECT 3.070 400.880 966.395 408.320 ;
        RECT 4.400 399.480 966.395 400.880 ;
        RECT 3.070 392.040 966.395 399.480 ;
        RECT 4.400 390.640 966.395 392.040 ;
        RECT 3.070 383.200 966.395 390.640 ;
        RECT 4.400 381.800 966.395 383.200 ;
        RECT 3.070 374.360 966.395 381.800 ;
        RECT 4.400 372.960 966.395 374.360 ;
        RECT 3.070 365.520 966.395 372.960 ;
        RECT 4.400 364.120 966.395 365.520 ;
        RECT 3.070 356.680 966.395 364.120 ;
        RECT 4.400 355.280 966.395 356.680 ;
        RECT 3.070 347.840 966.395 355.280 ;
        RECT 4.400 346.440 966.395 347.840 ;
        RECT 3.070 339.000 966.395 346.440 ;
        RECT 4.400 337.600 966.395 339.000 ;
        RECT 3.070 330.160 966.395 337.600 ;
        RECT 4.400 328.760 966.395 330.160 ;
        RECT 3.070 321.320 966.395 328.760 ;
        RECT 4.400 319.920 966.395 321.320 ;
        RECT 3.070 312.480 966.395 319.920 ;
        RECT 4.400 311.080 966.395 312.480 ;
        RECT 3.070 303.640 966.395 311.080 ;
        RECT 4.400 302.240 966.395 303.640 ;
        RECT 3.070 294.800 966.395 302.240 ;
        RECT 4.400 293.400 966.395 294.800 ;
        RECT 3.070 285.960 966.395 293.400 ;
        RECT 4.400 284.560 966.395 285.960 ;
        RECT 3.070 277.120 966.395 284.560 ;
        RECT 4.400 275.720 966.395 277.120 ;
        RECT 3.070 268.280 966.395 275.720 ;
        RECT 4.400 266.880 966.395 268.280 ;
        RECT 3.070 259.440 966.395 266.880 ;
        RECT 4.400 258.040 966.395 259.440 ;
        RECT 3.070 250.600 966.395 258.040 ;
        RECT 4.400 249.200 966.395 250.600 ;
        RECT 3.070 241.760 966.395 249.200 ;
        RECT 4.400 240.360 966.395 241.760 ;
        RECT 3.070 232.920 966.395 240.360 ;
        RECT 4.400 231.520 966.395 232.920 ;
        RECT 3.070 224.080 966.395 231.520 ;
        RECT 4.400 222.680 966.395 224.080 ;
        RECT 3.070 215.240 966.395 222.680 ;
        RECT 4.400 213.840 966.395 215.240 ;
        RECT 3.070 206.400 966.395 213.840 ;
        RECT 4.400 205.000 966.395 206.400 ;
        RECT 3.070 197.560 966.395 205.000 ;
        RECT 4.400 196.160 966.395 197.560 ;
        RECT 3.070 188.720 966.395 196.160 ;
        RECT 4.400 187.320 966.395 188.720 ;
        RECT 3.070 179.880 966.395 187.320 ;
        RECT 4.400 178.480 966.395 179.880 ;
        RECT 3.070 171.040 966.395 178.480 ;
        RECT 4.400 169.640 966.395 171.040 ;
        RECT 3.070 162.200 966.395 169.640 ;
        RECT 4.400 160.800 966.395 162.200 ;
        RECT 3.070 153.360 966.395 160.800 ;
        RECT 4.400 151.960 966.395 153.360 ;
        RECT 3.070 144.520 966.395 151.960 ;
        RECT 4.400 143.120 966.395 144.520 ;
        RECT 3.070 135.680 966.395 143.120 ;
        RECT 4.400 134.280 966.395 135.680 ;
        RECT 3.070 126.840 966.395 134.280 ;
        RECT 4.400 125.440 966.395 126.840 ;
        RECT 3.070 118.000 966.395 125.440 ;
        RECT 4.400 116.600 966.395 118.000 ;
        RECT 3.070 109.160 966.395 116.600 ;
        RECT 4.400 107.760 966.395 109.160 ;
        RECT 3.070 100.320 966.395 107.760 ;
        RECT 4.400 98.920 966.395 100.320 ;
        RECT 3.070 91.480 966.395 98.920 ;
        RECT 4.400 90.080 966.395 91.480 ;
        RECT 3.070 82.640 966.395 90.080 ;
        RECT 4.400 81.240 966.395 82.640 ;
        RECT 3.070 73.800 966.395 81.240 ;
        RECT 4.400 72.400 966.395 73.800 ;
        RECT 3.070 64.960 966.395 72.400 ;
        RECT 4.400 63.560 966.395 64.960 ;
        RECT 3.070 56.120 966.395 63.560 ;
        RECT 4.400 54.720 966.395 56.120 ;
        RECT 3.070 47.280 966.395 54.720 ;
        RECT 4.400 45.880 966.395 47.280 ;
        RECT 3.070 38.440 966.395 45.880 ;
        RECT 4.400 37.040 966.395 38.440 ;
        RECT 3.070 29.600 966.395 37.040 ;
        RECT 4.400 28.200 966.395 29.600 ;
        RECT 3.070 20.760 966.395 28.200 ;
        RECT 4.400 19.360 966.395 20.760 ;
        RECT 3.070 1.535 966.395 19.360 ;
      LAYER met4 ;
        RECT 63.775 10.240 97.440 313.985 ;
        RECT 99.840 10.240 174.240 313.985 ;
        RECT 176.640 10.240 251.040 313.985 ;
        RECT 253.440 10.240 327.840 313.985 ;
        RECT 330.240 10.240 404.640 313.985 ;
        RECT 407.040 10.240 481.440 313.985 ;
        RECT 483.840 10.240 558.240 313.985 ;
        RECT 560.640 10.240 635.040 313.985 ;
        RECT 637.440 10.240 651.985 313.985 ;
        RECT 63.775 1.535 651.985 10.240 ;
  END
END GPR
END LIBRARY

