module WBExecute (
  input      [31:0]   src0,
  input      [31:0]   src1,
  input      [31:0]   src2,
  input      [31:0]   src3,
  input      [31:0]   src4,
  input      [31:0]   src5,
  input      [5:0]    sel,
  input      [2:0]    zom,
  output reg [31:0]   result
);
endmodule