module REG32 (
  output     [31:0]   q,
  input               we,
  input      [31:0]   d,
  input               clk,
  input               reset
);
endmodule