module MUL16_U (
  input      [15:0]   src1,
  input      [15:0]   src2,
  output     [31:0]   result
);
endmodule