VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO MULADD_2
  CLASS BLOCK ;
  FOREIGN MULADD_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 100.000 ;
  PIN result[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END result[0]
  PIN result[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 4.000 ;
    END
  END result[10]
  PIN result[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 0.000 20.150 4.000 ;
    END
  END result[11]
  PIN result[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 4.000 ;
    END
  END result[12]
  PIN result[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END result[13]
  PIN result[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 4.000 ;
    END
  END result[14]
  PIN result[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 4.000 ;
    END
  END result[15]
  PIN result[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 4.000 ;
    END
  END result[16]
  PIN result[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 0.000 28.430 4.000 ;
    END
  END result[17]
  PIN result[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 4.000 ;
    END
  END result[18]
  PIN result[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 4.000 ;
    END
  END result[19]
  PIN result[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 0.000 6.350 4.000 ;
    END
  END result[1]
  PIN result[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END result[20]
  PIN result[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 4.000 ;
    END
  END result[21]
  PIN result[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END result[22]
  PIN result[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 4.000 ;
    END
  END result[23]
  PIN result[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 4.000 ;
    END
  END result[24]
  PIN result[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 4.000 ;
    END
  END result[25]
  PIN result[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END result[26]
  PIN result[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END result[27]
  PIN result[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END result[28]
  PIN result[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 0.000 44.990 4.000 ;
    END
  END result[29]
  PIN result[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END result[2]
  PIN result[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 0.000 46.370 4.000 ;
    END
  END result[30]
  PIN result[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 0.000 47.750 4.000 ;
    END
  END result[31]
  PIN result[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END result[32]
  PIN result[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 0.000 50.510 4.000 ;
    END
  END result[33]
  PIN result[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END result[34]
  PIN result[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 4.000 ;
    END
  END result[35]
  PIN result[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 0.000 54.650 4.000 ;
    END
  END result[36]
  PIN result[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END result[37]
  PIN result[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 0.000 57.410 4.000 ;
    END
  END result[38]
  PIN result[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 4.000 ;
    END
  END result[39]
  PIN result[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 0.000 9.110 4.000 ;
    END
  END result[3]
  PIN result[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END result[40]
  PIN result[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END result[41]
  PIN result[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END result[42]
  PIN result[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 4.000 ;
    END
  END result[43]
  PIN result[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 4.000 ;
    END
  END result[44]
  PIN result[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 0.000 67.070 4.000 ;
    END
  END result[45]
  PIN result[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 4.000 ;
    END
  END result[46]
  PIN result[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 4.000 ;
    END
  END result[47]
  PIN result[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END result[48]
  PIN result[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END result[49]
  PIN result[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 4.000 ;
    END
  END result[4]
  PIN result[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END result[50]
  PIN result[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 0.000 75.350 4.000 ;
    END
  END result[51]
  PIN result[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 4.000 ;
    END
  END result[52]
  PIN result[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 0.000 78.110 4.000 ;
    END
  END result[53]
  PIN result[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END result[54]
  PIN result[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END result[55]
  PIN result[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 4.000 ;
    END
  END result[56]
  PIN result[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 4.000 ;
    END
  END result[57]
  PIN result[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 4.000 ;
    END
  END result[58]
  PIN result[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 0.000 86.390 4.000 ;
    END
  END result[59]
  PIN result[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END result[5]
  PIN result[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END result[60]
  PIN result[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 0.000 89.150 4.000 ;
    END
  END result[61]
  PIN result[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END result[62]
  PIN result[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 0.000 91.910 4.000 ;
    END
  END result[63]
  PIN result[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END result[64]
  PIN result[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 4.000 ;
    END
  END result[65]
  PIN result[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END result[6]
  PIN result[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 0.000 14.630 4.000 ;
    END
  END result[7]
  PIN result[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 0.000 16.010 4.000 ;
    END
  END result[8]
  PIN result[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 0.000 17.390 4.000 ;
    END
  END result[9]
  PIN src1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 96.000 10.950 100.000 ;
    END
  END src1[0]
  PIN src1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 96.000 20.150 100.000 ;
    END
  END src1[10]
  PIN src1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 96.000 21.070 100.000 ;
    END
  END src1[11]
  PIN src1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 96.000 21.990 100.000 ;
    END
  END src1[12]
  PIN src1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 96.000 22.910 100.000 ;
    END
  END src1[13]
  PIN src1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 96.000 23.830 100.000 ;
    END
  END src1[14]
  PIN src1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 96.000 24.750 100.000 ;
    END
  END src1[15]
  PIN src1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 96.000 25.670 100.000 ;
    END
  END src1[16]
  PIN src1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 96.000 26.590 100.000 ;
    END
  END src1[17]
  PIN src1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 96.000 27.510 100.000 ;
    END
  END src1[18]
  PIN src1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 96.000 28.430 100.000 ;
    END
  END src1[19]
  PIN src1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 96.000 11.870 100.000 ;
    END
  END src1[1]
  PIN src1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 96.000 29.350 100.000 ;
    END
  END src1[20]
  PIN src1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 96.000 30.270 100.000 ;
    END
  END src1[21]
  PIN src1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 96.000 31.190 100.000 ;
    END
  END src1[22]
  PIN src1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 96.000 32.110 100.000 ;
    END
  END src1[23]
  PIN src1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.750 96.000 33.030 100.000 ;
    END
  END src1[24]
  PIN src1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 96.000 33.950 100.000 ;
    END
  END src1[25]
  PIN src1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 96.000 34.870 100.000 ;
    END
  END src1[26]
  PIN src1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 96.000 35.790 100.000 ;
    END
  END src1[27]
  PIN src1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 96.000 36.710 100.000 ;
    END
  END src1[28]
  PIN src1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 96.000 37.630 100.000 ;
    END
  END src1[29]
  PIN src1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 96.000 12.790 100.000 ;
    END
  END src1[2]
  PIN src1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 96.000 38.550 100.000 ;
    END
  END src1[30]
  PIN src1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 96.000 39.470 100.000 ;
    END
  END src1[31]
  PIN src1[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 96.000 40.390 100.000 ;
    END
  END src1[32]
  PIN src1[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 96.000 41.310 100.000 ;
    END
  END src1[33]
  PIN src1[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 96.000 42.230 100.000 ;
    END
  END src1[34]
  PIN src1[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 96.000 43.150 100.000 ;
    END
  END src1[35]
  PIN src1[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 96.000 44.070 100.000 ;
    END
  END src1[36]
  PIN src1[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 96.000 44.990 100.000 ;
    END
  END src1[37]
  PIN src1[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 96.000 45.910 100.000 ;
    END
  END src1[38]
  PIN src1[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 96.000 46.830 100.000 ;
    END
  END src1[39]
  PIN src1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.430 96.000 13.710 100.000 ;
    END
  END src1[3]
  PIN src1[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 96.000 47.750 100.000 ;
    END
  END src1[40]
  PIN src1[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 96.000 48.670 100.000 ;
    END
  END src1[41]
  PIN src1[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 96.000 49.590 100.000 ;
    END
  END src1[42]
  PIN src1[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 96.000 50.510 100.000 ;
    END
  END src1[43]
  PIN src1[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 96.000 51.430 100.000 ;
    END
  END src1[44]
  PIN src1[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 96.000 52.350 100.000 ;
    END
  END src1[45]
  PIN src1[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 96.000 53.270 100.000 ;
    END
  END src1[46]
  PIN src1[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 96.000 54.190 100.000 ;
    END
  END src1[47]
  PIN src1[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 96.000 55.110 100.000 ;
    END
  END src1[48]
  PIN src1[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 96.000 56.030 100.000 ;
    END
  END src1[49]
  PIN src1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 96.000 14.630 100.000 ;
    END
  END src1[4]
  PIN src1[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 96.000 56.950 100.000 ;
    END
  END src1[50]
  PIN src1[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 96.000 57.870 100.000 ;
    END
  END src1[51]
  PIN src1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 96.000 15.550 100.000 ;
    END
  END src1[5]
  PIN src1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 96.000 16.470 100.000 ;
    END
  END src1[6]
  PIN src1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 96.000 17.390 100.000 ;
    END
  END src1[7]
  PIN src1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 96.000 18.310 100.000 ;
    END
  END src1[8]
  PIN src1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 96.000 19.230 100.000 ;
    END
  END src1[9]
  PIN src2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 96.000 58.790 100.000 ;
    END
  END src2[0]
  PIN src2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 96.000 67.990 100.000 ;
    END
  END src2[10]
  PIN src2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 96.000 68.910 100.000 ;
    END
  END src2[11]
  PIN src2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 96.000 69.830 100.000 ;
    END
  END src2[12]
  PIN src2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 96.000 70.750 100.000 ;
    END
  END src2[13]
  PIN src2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 96.000 71.670 100.000 ;
    END
  END src2[14]
  PIN src2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 96.000 72.590 100.000 ;
    END
  END src2[15]
  PIN src2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 96.000 73.510 100.000 ;
    END
  END src2[16]
  PIN src2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 96.000 74.430 100.000 ;
    END
  END src2[17]
  PIN src2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 96.000 75.350 100.000 ;
    END
  END src2[18]
  PIN src2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 96.000 76.270 100.000 ;
    END
  END src2[19]
  PIN src2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 96.000 59.710 100.000 ;
    END
  END src2[1]
  PIN src2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 96.000 77.190 100.000 ;
    END
  END src2[20]
  PIN src2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 96.000 78.110 100.000 ;
    END
  END src2[21]
  PIN src2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 96.000 79.030 100.000 ;
    END
  END src2[22]
  PIN src2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 96.000 79.950 100.000 ;
    END
  END src2[23]
  PIN src2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 96.000 80.870 100.000 ;
    END
  END src2[24]
  PIN src2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 96.000 81.790 100.000 ;
    END
  END src2[25]
  PIN src2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 96.000 82.710 100.000 ;
    END
  END src2[26]
  PIN src2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 96.000 83.630 100.000 ;
    END
  END src2[27]
  PIN src2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 96.000 84.550 100.000 ;
    END
  END src2[28]
  PIN src2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 96.000 85.470 100.000 ;
    END
  END src2[29]
  PIN src2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 96.000 60.630 100.000 ;
    END
  END src2[2]
  PIN src2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 96.000 86.390 100.000 ;
    END
  END src2[30]
  PIN src2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 96.000 87.310 100.000 ;
    END
  END src2[31]
  PIN src2[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 96.000 88.230 100.000 ;
    END
  END src2[32]
  PIN src2[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 96.000 89.150 100.000 ;
    END
  END src2[33]
  PIN src2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 96.000 61.550 100.000 ;
    END
  END src2[3]
  PIN src2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 96.000 62.470 100.000 ;
    END
  END src2[4]
  PIN src2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 96.000 63.390 100.000 ;
    END
  END src2[5]
  PIN src2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 96.000 64.310 100.000 ;
    END
  END src2[6]
  PIN src2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 96.000 65.230 100.000 ;
    END
  END src2[7]
  PIN src2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 96.000 66.150 100.000 ;
    END
  END src2[8]
  PIN src2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 96.000 67.070 100.000 ;
    END
  END src2[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 15.840 10.640 17.440 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.080 10.640 39.680 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 60.320 10.640 61.920 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 82.560 10.640 84.160 87.280 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 26.960 10.640 28.560 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 49.200 10.640 50.800 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 71.440 10.640 73.040 87.280 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 94.300 87.125 ;
      LAYER met1 ;
        RECT 4.670 5.480 94.690 89.720 ;
      LAYER met2 ;
        RECT 4.700 95.720 10.390 96.000 ;
        RECT 11.230 95.720 11.310 96.000 ;
        RECT 12.150 95.720 12.230 96.000 ;
        RECT 13.070 95.720 13.150 96.000 ;
        RECT 13.990 95.720 14.070 96.000 ;
        RECT 14.910 95.720 14.990 96.000 ;
        RECT 15.830 95.720 15.910 96.000 ;
        RECT 16.750 95.720 16.830 96.000 ;
        RECT 17.670 95.720 17.750 96.000 ;
        RECT 18.590 95.720 18.670 96.000 ;
        RECT 19.510 95.720 19.590 96.000 ;
        RECT 20.430 95.720 20.510 96.000 ;
        RECT 21.350 95.720 21.430 96.000 ;
        RECT 22.270 95.720 22.350 96.000 ;
        RECT 23.190 95.720 23.270 96.000 ;
        RECT 24.110 95.720 24.190 96.000 ;
        RECT 25.030 95.720 25.110 96.000 ;
        RECT 25.950 95.720 26.030 96.000 ;
        RECT 26.870 95.720 26.950 96.000 ;
        RECT 27.790 95.720 27.870 96.000 ;
        RECT 28.710 95.720 28.790 96.000 ;
        RECT 29.630 95.720 29.710 96.000 ;
        RECT 30.550 95.720 30.630 96.000 ;
        RECT 31.470 95.720 31.550 96.000 ;
        RECT 32.390 95.720 32.470 96.000 ;
        RECT 33.310 95.720 33.390 96.000 ;
        RECT 34.230 95.720 34.310 96.000 ;
        RECT 35.150 95.720 35.230 96.000 ;
        RECT 36.070 95.720 36.150 96.000 ;
        RECT 36.990 95.720 37.070 96.000 ;
        RECT 37.910 95.720 37.990 96.000 ;
        RECT 38.830 95.720 38.910 96.000 ;
        RECT 39.750 95.720 39.830 96.000 ;
        RECT 40.670 95.720 40.750 96.000 ;
        RECT 41.590 95.720 41.670 96.000 ;
        RECT 42.510 95.720 42.590 96.000 ;
        RECT 43.430 95.720 43.510 96.000 ;
        RECT 44.350 95.720 44.430 96.000 ;
        RECT 45.270 95.720 45.350 96.000 ;
        RECT 46.190 95.720 46.270 96.000 ;
        RECT 47.110 95.720 47.190 96.000 ;
        RECT 48.030 95.720 48.110 96.000 ;
        RECT 48.950 95.720 49.030 96.000 ;
        RECT 49.870 95.720 49.950 96.000 ;
        RECT 50.790 95.720 50.870 96.000 ;
        RECT 51.710 95.720 51.790 96.000 ;
        RECT 52.630 95.720 52.710 96.000 ;
        RECT 53.550 95.720 53.630 96.000 ;
        RECT 54.470 95.720 54.550 96.000 ;
        RECT 55.390 95.720 55.470 96.000 ;
        RECT 56.310 95.720 56.390 96.000 ;
        RECT 57.230 95.720 57.310 96.000 ;
        RECT 58.150 95.720 58.230 96.000 ;
        RECT 59.070 95.720 59.150 96.000 ;
        RECT 59.990 95.720 60.070 96.000 ;
        RECT 60.910 95.720 60.990 96.000 ;
        RECT 61.830 95.720 61.910 96.000 ;
        RECT 62.750 95.720 62.830 96.000 ;
        RECT 63.670 95.720 63.750 96.000 ;
        RECT 64.590 95.720 64.670 96.000 ;
        RECT 65.510 95.720 65.590 96.000 ;
        RECT 66.430 95.720 66.510 96.000 ;
        RECT 67.350 95.720 67.430 96.000 ;
        RECT 68.270 95.720 68.350 96.000 ;
        RECT 69.190 95.720 69.270 96.000 ;
        RECT 70.110 95.720 70.190 96.000 ;
        RECT 71.030 95.720 71.110 96.000 ;
        RECT 71.950 95.720 72.030 96.000 ;
        RECT 72.870 95.720 72.950 96.000 ;
        RECT 73.790 95.720 73.870 96.000 ;
        RECT 74.710 95.720 74.790 96.000 ;
        RECT 75.630 95.720 75.710 96.000 ;
        RECT 76.550 95.720 76.630 96.000 ;
        RECT 77.470 95.720 77.550 96.000 ;
        RECT 78.390 95.720 78.470 96.000 ;
        RECT 79.310 95.720 79.390 96.000 ;
        RECT 80.230 95.720 80.310 96.000 ;
        RECT 81.150 95.720 81.230 96.000 ;
        RECT 82.070 95.720 82.150 96.000 ;
        RECT 82.990 95.720 83.070 96.000 ;
        RECT 83.910 95.720 83.990 96.000 ;
        RECT 84.830 95.720 84.910 96.000 ;
        RECT 85.750 95.720 85.830 96.000 ;
        RECT 86.670 95.720 86.750 96.000 ;
        RECT 87.590 95.720 87.670 96.000 ;
        RECT 88.510 95.720 88.590 96.000 ;
        RECT 89.430 95.720 94.660 96.000 ;
        RECT 4.700 4.280 94.660 95.720 ;
        RECT 5.250 4.000 5.790 4.280 ;
        RECT 6.630 4.000 7.170 4.280 ;
        RECT 8.010 4.000 8.550 4.280 ;
        RECT 9.390 4.000 9.930 4.280 ;
        RECT 10.770 4.000 11.310 4.280 ;
        RECT 12.150 4.000 12.690 4.280 ;
        RECT 13.530 4.000 14.070 4.280 ;
        RECT 14.910 4.000 15.450 4.280 ;
        RECT 16.290 4.000 16.830 4.280 ;
        RECT 17.670 4.000 18.210 4.280 ;
        RECT 19.050 4.000 19.590 4.280 ;
        RECT 20.430 4.000 20.970 4.280 ;
        RECT 21.810 4.000 22.350 4.280 ;
        RECT 23.190 4.000 23.730 4.280 ;
        RECT 24.570 4.000 25.110 4.280 ;
        RECT 25.950 4.000 26.490 4.280 ;
        RECT 27.330 4.000 27.870 4.280 ;
        RECT 28.710 4.000 29.250 4.280 ;
        RECT 30.090 4.000 30.630 4.280 ;
        RECT 31.470 4.000 32.010 4.280 ;
        RECT 32.850 4.000 33.390 4.280 ;
        RECT 34.230 4.000 34.770 4.280 ;
        RECT 35.610 4.000 36.150 4.280 ;
        RECT 36.990 4.000 37.530 4.280 ;
        RECT 38.370 4.000 38.910 4.280 ;
        RECT 39.750 4.000 40.290 4.280 ;
        RECT 41.130 4.000 41.670 4.280 ;
        RECT 42.510 4.000 43.050 4.280 ;
        RECT 43.890 4.000 44.430 4.280 ;
        RECT 45.270 4.000 45.810 4.280 ;
        RECT 46.650 4.000 47.190 4.280 ;
        RECT 48.030 4.000 48.570 4.280 ;
        RECT 49.410 4.000 49.950 4.280 ;
        RECT 50.790 4.000 51.330 4.280 ;
        RECT 52.170 4.000 52.710 4.280 ;
        RECT 53.550 4.000 54.090 4.280 ;
        RECT 54.930 4.000 55.470 4.280 ;
        RECT 56.310 4.000 56.850 4.280 ;
        RECT 57.690 4.000 58.230 4.280 ;
        RECT 59.070 4.000 59.610 4.280 ;
        RECT 60.450 4.000 60.990 4.280 ;
        RECT 61.830 4.000 62.370 4.280 ;
        RECT 63.210 4.000 63.750 4.280 ;
        RECT 64.590 4.000 65.130 4.280 ;
        RECT 65.970 4.000 66.510 4.280 ;
        RECT 67.350 4.000 67.890 4.280 ;
        RECT 68.730 4.000 69.270 4.280 ;
        RECT 70.110 4.000 70.650 4.280 ;
        RECT 71.490 4.000 72.030 4.280 ;
        RECT 72.870 4.000 73.410 4.280 ;
        RECT 74.250 4.000 74.790 4.280 ;
        RECT 75.630 4.000 76.170 4.280 ;
        RECT 77.010 4.000 77.550 4.280 ;
        RECT 78.390 4.000 78.930 4.280 ;
        RECT 79.770 4.000 80.310 4.280 ;
        RECT 81.150 4.000 81.690 4.280 ;
        RECT 82.530 4.000 83.070 4.280 ;
        RECT 83.910 4.000 84.450 4.280 ;
        RECT 85.290 4.000 85.830 4.280 ;
        RECT 86.670 4.000 87.210 4.280 ;
        RECT 88.050 4.000 88.590 4.280 ;
        RECT 89.430 4.000 89.970 4.280 ;
        RECT 90.810 4.000 91.350 4.280 ;
        RECT 92.190 4.000 92.730 4.280 ;
        RECT 93.570 4.000 94.110 4.280 ;
      LAYER met3 ;
        RECT 12.945 10.715 87.795 87.205 ;
      LAYER met4 ;
        RECT 53.655 11.735 59.920 76.665 ;
        RECT 62.320 11.735 71.040 76.665 ;
        RECT 73.440 11.735 82.160 76.665 ;
        RECT 84.560 11.735 87.105 76.665 ;
  END
END MULADD_2
END LIBRARY

