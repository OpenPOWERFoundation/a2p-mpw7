module MUL17_S (
  input      [16:0]   src1,
  input      [16:0]   src2,
  output     [33:0]   result
);
endmodule