VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO InstructionCache
  CLASS BLOCK ;
  FOREIGN InstructionCache ;
  ORIGIN 0.000 0.000 ;
  SIZE 650.000 BY 250.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.530 246.000 627.810 250.000 ;
    END
  END clk
  PIN io_cpu_decode_cacheMiss
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 246.000 20.610 250.000 ;
    END
  END io_cpu_decode_cacheMiss
  PIN io_cpu_decode_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 246.000 56.490 250.000 ;
    END
  END io_cpu_decode_data[0]
  PIN io_cpu_decode_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.850 246.000 233.130 250.000 ;
    END
  END io_cpu_decode_data[10]
  PIN io_cpu_decode_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 246.000 248.310 250.000 ;
    END
  END io_cpu_decode_data[11]
  PIN io_cpu_decode_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.210 246.000 263.490 250.000 ;
    END
  END io_cpu_decode_data[12]
  PIN io_cpu_decode_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.390 246.000 278.670 250.000 ;
    END
  END io_cpu_decode_data[13]
  PIN io_cpu_decode_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 246.000 293.850 250.000 ;
    END
  END io_cpu_decode_data[14]
  PIN io_cpu_decode_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 246.000 309.030 250.000 ;
    END
  END io_cpu_decode_data[15]
  PIN io_cpu_decode_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.930 246.000 324.210 250.000 ;
    END
  END io_cpu_decode_data[16]
  PIN io_cpu_decode_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.110 246.000 339.390 250.000 ;
    END
  END io_cpu_decode_data[17]
  PIN io_cpu_decode_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 246.000 354.570 250.000 ;
    END
  END io_cpu_decode_data[18]
  PIN io_cpu_decode_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.470 246.000 369.750 250.000 ;
    END
  END io_cpu_decode_data[19]
  PIN io_cpu_decode_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 246.000 75.810 250.000 ;
    END
  END io_cpu_decode_data[1]
  PIN io_cpu_decode_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.650 246.000 384.930 250.000 ;
    END
  END io_cpu_decode_data[20]
  PIN io_cpu_decode_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.830 246.000 400.110 250.000 ;
    END
  END io_cpu_decode_data[21]
  PIN io_cpu_decode_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.010 246.000 415.290 250.000 ;
    END
  END io_cpu_decode_data[22]
  PIN io_cpu_decode_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.190 246.000 430.470 250.000 ;
    END
  END io_cpu_decode_data[23]
  PIN io_cpu_decode_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.370 246.000 445.650 250.000 ;
    END
  END io_cpu_decode_data[24]
  PIN io_cpu_decode_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 246.000 460.830 250.000 ;
    END
  END io_cpu_decode_data[25]
  PIN io_cpu_decode_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.730 246.000 476.010 250.000 ;
    END
  END io_cpu_decode_data[26]
  PIN io_cpu_decode_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.910 246.000 491.190 250.000 ;
    END
  END io_cpu_decode_data[27]
  PIN io_cpu_decode_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.090 246.000 506.370 250.000 ;
    END
  END io_cpu_decode_data[28]
  PIN io_cpu_decode_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.270 246.000 521.550 250.000 ;
    END
  END io_cpu_decode_data[29]
  PIN io_cpu_decode_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 246.000 95.130 250.000 ;
    END
  END io_cpu_decode_data[2]
  PIN io_cpu_decode_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.450 246.000 536.730 250.000 ;
    END
  END io_cpu_decode_data[30]
  PIN io_cpu_decode_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.630 246.000 551.910 250.000 ;
    END
  END io_cpu_decode_data[31]
  PIN io_cpu_decode_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 246.000 114.450 250.000 ;
    END
  END io_cpu_decode_data[3]
  PIN io_cpu_decode_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 246.000 133.770 250.000 ;
    END
  END io_cpu_decode_data[4]
  PIN io_cpu_decode_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 246.000 150.330 250.000 ;
    END
  END io_cpu_decode_data[5]
  PIN io_cpu_decode_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 246.000 166.890 250.000 ;
    END
  END io_cpu_decode_data[6]
  PIN io_cpu_decode_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.170 246.000 183.450 250.000 ;
    END
  END io_cpu_decode_data[7]
  PIN io_cpu_decode_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 246.000 200.010 250.000 ;
    END
  END io_cpu_decode_data[8]
  PIN io_cpu_decode_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 246.000 216.570 250.000 ;
    END
  END io_cpu_decode_data[9]
  PIN io_cpu_decode_error
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 246.000 21.990 250.000 ;
    END
  END io_cpu_decode_error
  PIN io_cpu_decode_exceptionType[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 246.000 57.870 250.000 ;
    END
  END io_cpu_decode_exceptionType[0]
  PIN io_cpu_decode_exceptionType[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 246.000 77.190 250.000 ;
    END
  END io_cpu_decode_exceptionType[1]
  PIN io_cpu_decode_exceptionType[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 246.000 96.510 250.000 ;
    END
  END io_cpu_decode_exceptionType[2]
  PIN io_cpu_decode_exceptionType[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 246.000 115.830 250.000 ;
    END
  END io_cpu_decode_exceptionType[3]
  PIN io_cpu_decode_isStuck
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 246.000 23.370 250.000 ;
    END
  END io_cpu_decode_isStuck
  PIN io_cpu_decode_isUser
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 246.000 24.750 250.000 ;
    END
  END io_cpu_decode_isUser
  PIN io_cpu_decode_isValid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 246.000 26.130 250.000 ;
    END
  END io_cpu_decode_isValid
  PIN io_cpu_decode_mmuException
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 246.000 27.510 250.000 ;
    END
  END io_cpu_decode_mmuException
  PIN io_cpu_decode_mmuRefilling
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 246.000 28.890 250.000 ;
    END
  END io_cpu_decode_mmuRefilling
  PIN io_cpu_decode_pc[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 246.000 59.250 250.000 ;
    END
  END io_cpu_decode_pc[0]
  PIN io_cpu_decode_pc[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.230 246.000 234.510 250.000 ;
    END
  END io_cpu_decode_pc[10]
  PIN io_cpu_decode_pc[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 246.000 249.690 250.000 ;
    END
  END io_cpu_decode_pc[11]
  PIN io_cpu_decode_pc[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 246.000 264.870 250.000 ;
    END
  END io_cpu_decode_pc[12]
  PIN io_cpu_decode_pc[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 246.000 280.050 250.000 ;
    END
  END io_cpu_decode_pc[13]
  PIN io_cpu_decode_pc[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 246.000 295.230 250.000 ;
    END
  END io_cpu_decode_pc[14]
  PIN io_cpu_decode_pc[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.130 246.000 310.410 250.000 ;
    END
  END io_cpu_decode_pc[15]
  PIN io_cpu_decode_pc[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 246.000 325.590 250.000 ;
    END
  END io_cpu_decode_pc[16]
  PIN io_cpu_decode_pc[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.490 246.000 340.770 250.000 ;
    END
  END io_cpu_decode_pc[17]
  PIN io_cpu_decode_pc[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.670 246.000 355.950 250.000 ;
    END
  END io_cpu_decode_pc[18]
  PIN io_cpu_decode_pc[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.850 246.000 371.130 250.000 ;
    END
  END io_cpu_decode_pc[19]
  PIN io_cpu_decode_pc[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 246.000 78.570 250.000 ;
    END
  END io_cpu_decode_pc[1]
  PIN io_cpu_decode_pc[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.030 246.000 386.310 250.000 ;
    END
  END io_cpu_decode_pc[20]
  PIN io_cpu_decode_pc[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.210 246.000 401.490 250.000 ;
    END
  END io_cpu_decode_pc[21]
  PIN io_cpu_decode_pc[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.390 246.000 416.670 250.000 ;
    END
  END io_cpu_decode_pc[22]
  PIN io_cpu_decode_pc[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 246.000 431.850 250.000 ;
    END
  END io_cpu_decode_pc[23]
  PIN io_cpu_decode_pc[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.750 246.000 447.030 250.000 ;
    END
  END io_cpu_decode_pc[24]
  PIN io_cpu_decode_pc[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.930 246.000 462.210 250.000 ;
    END
  END io_cpu_decode_pc[25]
  PIN io_cpu_decode_pc[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.110 246.000 477.390 250.000 ;
    END
  END io_cpu_decode_pc[26]
  PIN io_cpu_decode_pc[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.290 246.000 492.570 250.000 ;
    END
  END io_cpu_decode_pc[27]
  PIN io_cpu_decode_pc[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.470 246.000 507.750 250.000 ;
    END
  END io_cpu_decode_pc[28]
  PIN io_cpu_decode_pc[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.650 246.000 522.930 250.000 ;
    END
  END io_cpu_decode_pc[29]
  PIN io_cpu_decode_pc[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 246.000 97.890 250.000 ;
    END
  END io_cpu_decode_pc[2]
  PIN io_cpu_decode_pc[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 246.000 538.110 250.000 ;
    END
  END io_cpu_decode_pc[30]
  PIN io_cpu_decode_pc[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.010 246.000 553.290 250.000 ;
    END
  END io_cpu_decode_pc[31]
  PIN io_cpu_decode_pc[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 246.000 117.210 250.000 ;
    END
  END io_cpu_decode_pc[3]
  PIN io_cpu_decode_pc[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.870 246.000 135.150 250.000 ;
    END
  END io_cpu_decode_pc[4]
  PIN io_cpu_decode_pc[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 246.000 151.710 250.000 ;
    END
  END io_cpu_decode_pc[5]
  PIN io_cpu_decode_pc[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 246.000 168.270 250.000 ;
    END
  END io_cpu_decode_pc[6]
  PIN io_cpu_decode_pc[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.550 246.000 184.830 250.000 ;
    END
  END io_cpu_decode_pc[7]
  PIN io_cpu_decode_pc[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.110 246.000 201.390 250.000 ;
    END
  END io_cpu_decode_pc[8]
  PIN io_cpu_decode_pc[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 246.000 217.950 250.000 ;
    END
  END io_cpu_decode_pc[9]
  PIN io_cpu_decode_physicalAddress[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 246.000 60.630 250.000 ;
    END
  END io_cpu_decode_physicalAddress[0]
  PIN io_cpu_decode_physicalAddress[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.610 246.000 235.890 250.000 ;
    END
  END io_cpu_decode_physicalAddress[10]
  PIN io_cpu_decode_physicalAddress[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.790 246.000 251.070 250.000 ;
    END
  END io_cpu_decode_physicalAddress[11]
  PIN io_cpu_decode_physicalAddress[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.970 246.000 266.250 250.000 ;
    END
  END io_cpu_decode_physicalAddress[12]
  PIN io_cpu_decode_physicalAddress[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 246.000 281.430 250.000 ;
    END
  END io_cpu_decode_physicalAddress[13]
  PIN io_cpu_decode_physicalAddress[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 246.000 296.610 250.000 ;
    END
  END io_cpu_decode_physicalAddress[14]
  PIN io_cpu_decode_physicalAddress[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.510 246.000 311.790 250.000 ;
    END
  END io_cpu_decode_physicalAddress[15]
  PIN io_cpu_decode_physicalAddress[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 246.000 326.970 250.000 ;
    END
  END io_cpu_decode_physicalAddress[16]
  PIN io_cpu_decode_physicalAddress[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.870 246.000 342.150 250.000 ;
    END
  END io_cpu_decode_physicalAddress[17]
  PIN io_cpu_decode_physicalAddress[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 246.000 357.330 250.000 ;
    END
  END io_cpu_decode_physicalAddress[18]
  PIN io_cpu_decode_physicalAddress[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.230 246.000 372.510 250.000 ;
    END
  END io_cpu_decode_physicalAddress[19]
  PIN io_cpu_decode_physicalAddress[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 246.000 79.950 250.000 ;
    END
  END io_cpu_decode_physicalAddress[1]
  PIN io_cpu_decode_physicalAddress[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.410 246.000 387.690 250.000 ;
    END
  END io_cpu_decode_physicalAddress[20]
  PIN io_cpu_decode_physicalAddress[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 246.000 402.870 250.000 ;
    END
  END io_cpu_decode_physicalAddress[21]
  PIN io_cpu_decode_physicalAddress[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.770 246.000 418.050 250.000 ;
    END
  END io_cpu_decode_physicalAddress[22]
  PIN io_cpu_decode_physicalAddress[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.950 246.000 433.230 250.000 ;
    END
  END io_cpu_decode_physicalAddress[23]
  PIN io_cpu_decode_physicalAddress[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.130 246.000 448.410 250.000 ;
    END
  END io_cpu_decode_physicalAddress[24]
  PIN io_cpu_decode_physicalAddress[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.310 246.000 463.590 250.000 ;
    END
  END io_cpu_decode_physicalAddress[25]
  PIN io_cpu_decode_physicalAddress[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.490 246.000 478.770 250.000 ;
    END
  END io_cpu_decode_physicalAddress[26]
  PIN io_cpu_decode_physicalAddress[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.670 246.000 493.950 250.000 ;
    END
  END io_cpu_decode_physicalAddress[27]
  PIN io_cpu_decode_physicalAddress[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 246.000 509.130 250.000 ;
    END
  END io_cpu_decode_physicalAddress[28]
  PIN io_cpu_decode_physicalAddress[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.030 246.000 524.310 250.000 ;
    END
  END io_cpu_decode_physicalAddress[29]
  PIN io_cpu_decode_physicalAddress[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 246.000 99.270 250.000 ;
    END
  END io_cpu_decode_physicalAddress[2]
  PIN io_cpu_decode_physicalAddress[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.210 246.000 539.490 250.000 ;
    END
  END io_cpu_decode_physicalAddress[30]
  PIN io_cpu_decode_physicalAddress[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.390 246.000 554.670 250.000 ;
    END
  END io_cpu_decode_physicalAddress[31]
  PIN io_cpu_decode_physicalAddress[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.310 246.000 118.590 250.000 ;
    END
  END io_cpu_decode_physicalAddress[3]
  PIN io_cpu_decode_physicalAddress[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.250 246.000 136.530 250.000 ;
    END
  END io_cpu_decode_physicalAddress[4]
  PIN io_cpu_decode_physicalAddress[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 246.000 153.090 250.000 ;
    END
  END io_cpu_decode_physicalAddress[5]
  PIN io_cpu_decode_physicalAddress[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 246.000 169.650 250.000 ;
    END
  END io_cpu_decode_physicalAddress[6]
  PIN io_cpu_decode_physicalAddress[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 246.000 186.210 250.000 ;
    END
  END io_cpu_decode_physicalAddress[7]
  PIN io_cpu_decode_physicalAddress[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.490 246.000 202.770 250.000 ;
    END
  END io_cpu_decode_physicalAddress[8]
  PIN io_cpu_decode_physicalAddress[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 246.000 219.330 250.000 ;
    END
  END io_cpu_decode_physicalAddress[9]
  PIN io_cpu_fetch_bypassTranslation
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 246.000 30.270 250.000 ;
    END
  END io_cpu_fetch_bypassTranslation
  PIN io_cpu_fetch_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 246.000 62.010 250.000 ;
    END
  END io_cpu_fetch_data[0]
  PIN io_cpu_fetch_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.990 246.000 237.270 250.000 ;
    END
  END io_cpu_fetch_data[10]
  PIN io_cpu_fetch_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 246.000 252.450 250.000 ;
    END
  END io_cpu_fetch_data[11]
  PIN io_cpu_fetch_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 246.000 267.630 250.000 ;
    END
  END io_cpu_fetch_data[12]
  PIN io_cpu_fetch_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.530 246.000 282.810 250.000 ;
    END
  END io_cpu_fetch_data[13]
  PIN io_cpu_fetch_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.710 246.000 297.990 250.000 ;
    END
  END io_cpu_fetch_data[14]
  PIN io_cpu_fetch_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 246.000 313.170 250.000 ;
    END
  END io_cpu_fetch_data[15]
  PIN io_cpu_fetch_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.070 246.000 328.350 250.000 ;
    END
  END io_cpu_fetch_data[16]
  PIN io_cpu_fetch_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.250 246.000 343.530 250.000 ;
    END
  END io_cpu_fetch_data[17]
  PIN io_cpu_fetch_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.430 246.000 358.710 250.000 ;
    END
  END io_cpu_fetch_data[18]
  PIN io_cpu_fetch_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 246.000 373.890 250.000 ;
    END
  END io_cpu_fetch_data[19]
  PIN io_cpu_fetch_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 246.000 81.330 250.000 ;
    END
  END io_cpu_fetch_data[1]
  PIN io_cpu_fetch_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.790 246.000 389.070 250.000 ;
    END
  END io_cpu_fetch_data[20]
  PIN io_cpu_fetch_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.970 246.000 404.250 250.000 ;
    END
  END io_cpu_fetch_data[21]
  PIN io_cpu_fetch_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.150 246.000 419.430 250.000 ;
    END
  END io_cpu_fetch_data[22]
  PIN io_cpu_fetch_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.330 246.000 434.610 250.000 ;
    END
  END io_cpu_fetch_data[23]
  PIN io_cpu_fetch_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 246.000 449.790 250.000 ;
    END
  END io_cpu_fetch_data[24]
  PIN io_cpu_fetch_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.690 246.000 464.970 250.000 ;
    END
  END io_cpu_fetch_data[25]
  PIN io_cpu_fetch_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 246.000 480.150 250.000 ;
    END
  END io_cpu_fetch_data[26]
  PIN io_cpu_fetch_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.050 246.000 495.330 250.000 ;
    END
  END io_cpu_fetch_data[27]
  PIN io_cpu_fetch_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.230 246.000 510.510 250.000 ;
    END
  END io_cpu_fetch_data[28]
  PIN io_cpu_fetch_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.410 246.000 525.690 250.000 ;
    END
  END io_cpu_fetch_data[29]
  PIN io_cpu_fetch_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 246.000 100.650 250.000 ;
    END
  END io_cpu_fetch_data[2]
  PIN io_cpu_fetch_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.590 246.000 540.870 250.000 ;
    END
  END io_cpu_fetch_data[30]
  PIN io_cpu_fetch_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.770 246.000 556.050 250.000 ;
    END
  END io_cpu_fetch_data[31]
  PIN io_cpu_fetch_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 246.000 119.970 250.000 ;
    END
  END io_cpu_fetch_data[3]
  PIN io_cpu_fetch_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 246.000 137.910 250.000 ;
    END
  END io_cpu_fetch_data[4]
  PIN io_cpu_fetch_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.190 246.000 154.470 250.000 ;
    END
  END io_cpu_fetch_data[5]
  PIN io_cpu_fetch_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 246.000 171.030 250.000 ;
    END
  END io_cpu_fetch_data[6]
  PIN io_cpu_fetch_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 246.000 187.590 250.000 ;
    END
  END io_cpu_fetch_data[7]
  PIN io_cpu_fetch_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.870 246.000 204.150 250.000 ;
    END
  END io_cpu_fetch_data[8]
  PIN io_cpu_fetch_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.430 246.000 220.710 250.000 ;
    END
  END io_cpu_fetch_data[9]
  PIN io_cpu_fetch_exceptionType[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 246.000 63.390 250.000 ;
    END
  END io_cpu_fetch_exceptionType[0]
  PIN io_cpu_fetch_exceptionType[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 246.000 82.710 250.000 ;
    END
  END io_cpu_fetch_exceptionType[1]
  PIN io_cpu_fetch_exceptionType[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.750 246.000 102.030 250.000 ;
    END
  END io_cpu_fetch_exceptionType[2]
  PIN io_cpu_fetch_exceptionType[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.070 246.000 121.350 250.000 ;
    END
  END io_cpu_fetch_exceptionType[3]
  PIN io_cpu_fetch_haltIt
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 246.000 31.650 250.000 ;
    END
  END io_cpu_fetch_haltIt
  PIN io_cpu_fetch_isRemoved
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.750 246.000 33.030 250.000 ;
    END
  END io_cpu_fetch_isRemoved
  PIN io_cpu_fetch_isStuck
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.130 246.000 34.410 250.000 ;
    END
  END io_cpu_fetch_isStuck
  PIN io_cpu_fetch_isValid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 246.000 35.790 250.000 ;
    END
  END io_cpu_fetch_isValid
  PIN io_cpu_fetch_mmuBus_busy
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 246.000 37.170 250.000 ;
    END
  END io_cpu_fetch_mmuBus_busy
  PIN io_cpu_fetch_mmuBus_cmd_bypassTranslation
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 246.000 38.550 250.000 ;
    END
  END io_cpu_fetch_mmuBus_cmd_bypassTranslation
  PIN io_cpu_fetch_mmuBus_cmd_isValid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 246.000 39.930 250.000 ;
    END
  END io_cpu_fetch_mmuBus_cmd_isValid
  PIN io_cpu_fetch_mmuBus_cmd_virtualAddress[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 246.000 64.770 250.000 ;
    END
  END io_cpu_fetch_mmuBus_cmd_virtualAddress[0]
  PIN io_cpu_fetch_mmuBus_cmd_virtualAddress[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 246.000 238.650 250.000 ;
    END
  END io_cpu_fetch_mmuBus_cmd_virtualAddress[10]
  PIN io_cpu_fetch_mmuBus_cmd_virtualAddress[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.550 246.000 253.830 250.000 ;
    END
  END io_cpu_fetch_mmuBus_cmd_virtualAddress[11]
  PIN io_cpu_fetch_mmuBus_cmd_virtualAddress[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.730 246.000 269.010 250.000 ;
    END
  END io_cpu_fetch_mmuBus_cmd_virtualAddress[12]
  PIN io_cpu_fetch_mmuBus_cmd_virtualAddress[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.910 246.000 284.190 250.000 ;
    END
  END io_cpu_fetch_mmuBus_cmd_virtualAddress[13]
  PIN io_cpu_fetch_mmuBus_cmd_virtualAddress[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.090 246.000 299.370 250.000 ;
    END
  END io_cpu_fetch_mmuBus_cmd_virtualAddress[14]
  PIN io_cpu_fetch_mmuBus_cmd_virtualAddress[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.270 246.000 314.550 250.000 ;
    END
  END io_cpu_fetch_mmuBus_cmd_virtualAddress[15]
  PIN io_cpu_fetch_mmuBus_cmd_virtualAddress[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.450 246.000 329.730 250.000 ;
    END
  END io_cpu_fetch_mmuBus_cmd_virtualAddress[16]
  PIN io_cpu_fetch_mmuBus_cmd_virtualAddress[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 246.000 344.910 250.000 ;
    END
  END io_cpu_fetch_mmuBus_cmd_virtualAddress[17]
  PIN io_cpu_fetch_mmuBus_cmd_virtualAddress[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.810 246.000 360.090 250.000 ;
    END
  END io_cpu_fetch_mmuBus_cmd_virtualAddress[18]
  PIN io_cpu_fetch_mmuBus_cmd_virtualAddress[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.990 246.000 375.270 250.000 ;
    END
  END io_cpu_fetch_mmuBus_cmd_virtualAddress[19]
  PIN io_cpu_fetch_mmuBus_cmd_virtualAddress[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 246.000 84.090 250.000 ;
    END
  END io_cpu_fetch_mmuBus_cmd_virtualAddress[1]
  PIN io_cpu_fetch_mmuBus_cmd_virtualAddress[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.170 246.000 390.450 250.000 ;
    END
  END io_cpu_fetch_mmuBus_cmd_virtualAddress[20]
  PIN io_cpu_fetch_mmuBus_cmd_virtualAddress[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.350 246.000 405.630 250.000 ;
    END
  END io_cpu_fetch_mmuBus_cmd_virtualAddress[21]
  PIN io_cpu_fetch_mmuBus_cmd_virtualAddress[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.530 246.000 420.810 250.000 ;
    END
  END io_cpu_fetch_mmuBus_cmd_virtualAddress[22]
  PIN io_cpu_fetch_mmuBus_cmd_virtualAddress[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.710 246.000 435.990 250.000 ;
    END
  END io_cpu_fetch_mmuBus_cmd_virtualAddress[23]
  PIN io_cpu_fetch_mmuBus_cmd_virtualAddress[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 246.000 451.170 250.000 ;
    END
  END io_cpu_fetch_mmuBus_cmd_virtualAddress[24]
  PIN io_cpu_fetch_mmuBus_cmd_virtualAddress[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.070 246.000 466.350 250.000 ;
    END
  END io_cpu_fetch_mmuBus_cmd_virtualAddress[25]
  PIN io_cpu_fetch_mmuBus_cmd_virtualAddress[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.250 246.000 481.530 250.000 ;
    END
  END io_cpu_fetch_mmuBus_cmd_virtualAddress[26]
  PIN io_cpu_fetch_mmuBus_cmd_virtualAddress[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.430 246.000 496.710 250.000 ;
    END
  END io_cpu_fetch_mmuBus_cmd_virtualAddress[27]
  PIN io_cpu_fetch_mmuBus_cmd_virtualAddress[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.610 246.000 511.890 250.000 ;
    END
  END io_cpu_fetch_mmuBus_cmd_virtualAddress[28]
  PIN io_cpu_fetch_mmuBus_cmd_virtualAddress[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.790 246.000 527.070 250.000 ;
    END
  END io_cpu_fetch_mmuBus_cmd_virtualAddress[29]
  PIN io_cpu_fetch_mmuBus_cmd_virtualAddress[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 246.000 103.410 250.000 ;
    END
  END io_cpu_fetch_mmuBus_cmd_virtualAddress[2]
  PIN io_cpu_fetch_mmuBus_cmd_virtualAddress[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.970 246.000 542.250 250.000 ;
    END
  END io_cpu_fetch_mmuBus_cmd_virtualAddress[30]
  PIN io_cpu_fetch_mmuBus_cmd_virtualAddress[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 246.000 557.430 250.000 ;
    END
  END io_cpu_fetch_mmuBus_cmd_virtualAddress[31]
  PIN io_cpu_fetch_mmuBus_cmd_virtualAddress[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 246.000 122.730 250.000 ;
    END
  END io_cpu_fetch_mmuBus_cmd_virtualAddress[3]
  PIN io_cpu_fetch_mmuBus_cmd_virtualAddress[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 246.000 139.290 250.000 ;
    END
  END io_cpu_fetch_mmuBus_cmd_virtualAddress[4]
  PIN io_cpu_fetch_mmuBus_cmd_virtualAddress[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 246.000 155.850 250.000 ;
    END
  END io_cpu_fetch_mmuBus_cmd_virtualAddress[5]
  PIN io_cpu_fetch_mmuBus_cmd_virtualAddress[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.130 246.000 172.410 250.000 ;
    END
  END io_cpu_fetch_mmuBus_cmd_virtualAddress[6]
  PIN io_cpu_fetch_mmuBus_cmd_virtualAddress[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.690 246.000 188.970 250.000 ;
    END
  END io_cpu_fetch_mmuBus_cmd_virtualAddress[7]
  PIN io_cpu_fetch_mmuBus_cmd_virtualAddress[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 246.000 205.530 250.000 ;
    END
  END io_cpu_fetch_mmuBus_cmd_virtualAddress[8]
  PIN io_cpu_fetch_mmuBus_cmd_virtualAddress[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.810 246.000 222.090 250.000 ;
    END
  END io_cpu_fetch_mmuBus_cmd_virtualAddress[9]
  PIN io_cpu_fetch_mmuBus_end
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 246.000 41.310 250.000 ;
    END
  END io_cpu_fetch_mmuBus_end
  PIN io_cpu_fetch_mmuBus_rsp_allowExecute
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 246.000 42.690 250.000 ;
    END
  END io_cpu_fetch_mmuBus_rsp_allowExecute
  PIN io_cpu_fetch_mmuBus_rsp_allowRead
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 246.000 44.070 250.000 ;
    END
  END io_cpu_fetch_mmuBus_rsp_allowRead
  PIN io_cpu_fetch_mmuBus_rsp_allowWrite
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 246.000 45.450 250.000 ;
    END
  END io_cpu_fetch_mmuBus_rsp_allowWrite
  PIN io_cpu_fetch_mmuBus_rsp_exception
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 246.000 46.830 250.000 ;
    END
  END io_cpu_fetch_mmuBus_rsp_exception
  PIN io_cpu_fetch_mmuBus_rsp_isIoAccess
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 246.000 48.210 250.000 ;
    END
  END io_cpu_fetch_mmuBus_rsp_isIoAccess
  PIN io_cpu_fetch_mmuBus_rsp_physicalAddress[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 246.000 66.150 250.000 ;
    END
  END io_cpu_fetch_mmuBus_rsp_physicalAddress[0]
  PIN io_cpu_fetch_mmuBus_rsp_physicalAddress[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.750 246.000 240.030 250.000 ;
    END
  END io_cpu_fetch_mmuBus_rsp_physicalAddress[10]
  PIN io_cpu_fetch_mmuBus_rsp_physicalAddress[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 246.000 255.210 250.000 ;
    END
  END io_cpu_fetch_mmuBus_rsp_physicalAddress[11]
  PIN io_cpu_fetch_mmuBus_rsp_physicalAddress[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 246.000 270.390 250.000 ;
    END
  END io_cpu_fetch_mmuBus_rsp_physicalAddress[12]
  PIN io_cpu_fetch_mmuBus_rsp_physicalAddress[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.290 246.000 285.570 250.000 ;
    END
  END io_cpu_fetch_mmuBus_rsp_physicalAddress[13]
  PIN io_cpu_fetch_mmuBus_rsp_physicalAddress[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.470 246.000 300.750 250.000 ;
    END
  END io_cpu_fetch_mmuBus_rsp_physicalAddress[14]
  PIN io_cpu_fetch_mmuBus_rsp_physicalAddress[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 246.000 315.930 250.000 ;
    END
  END io_cpu_fetch_mmuBus_rsp_physicalAddress[15]
  PIN io_cpu_fetch_mmuBus_rsp_physicalAddress[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 246.000 331.110 250.000 ;
    END
  END io_cpu_fetch_mmuBus_rsp_physicalAddress[16]
  PIN io_cpu_fetch_mmuBus_rsp_physicalAddress[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.010 246.000 346.290 250.000 ;
    END
  END io_cpu_fetch_mmuBus_rsp_physicalAddress[17]
  PIN io_cpu_fetch_mmuBus_rsp_physicalAddress[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.190 246.000 361.470 250.000 ;
    END
  END io_cpu_fetch_mmuBus_rsp_physicalAddress[18]
  PIN io_cpu_fetch_mmuBus_rsp_physicalAddress[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.370 246.000 376.650 250.000 ;
    END
  END io_cpu_fetch_mmuBus_rsp_physicalAddress[19]
  PIN io_cpu_fetch_mmuBus_rsp_physicalAddress[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 246.000 85.470 250.000 ;
    END
  END io_cpu_fetch_mmuBus_rsp_physicalAddress[1]
  PIN io_cpu_fetch_mmuBus_rsp_physicalAddress[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.550 246.000 391.830 250.000 ;
    END
  END io_cpu_fetch_mmuBus_rsp_physicalAddress[20]
  PIN io_cpu_fetch_mmuBus_rsp_physicalAddress[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.730 246.000 407.010 250.000 ;
    END
  END io_cpu_fetch_mmuBus_rsp_physicalAddress[21]
  PIN io_cpu_fetch_mmuBus_rsp_physicalAddress[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 246.000 422.190 250.000 ;
    END
  END io_cpu_fetch_mmuBus_rsp_physicalAddress[22]
  PIN io_cpu_fetch_mmuBus_rsp_physicalAddress[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.090 246.000 437.370 250.000 ;
    END
  END io_cpu_fetch_mmuBus_rsp_physicalAddress[23]
  PIN io_cpu_fetch_mmuBus_rsp_physicalAddress[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.270 246.000 452.550 250.000 ;
    END
  END io_cpu_fetch_mmuBus_rsp_physicalAddress[24]
  PIN io_cpu_fetch_mmuBus_rsp_physicalAddress[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.450 246.000 467.730 250.000 ;
    END
  END io_cpu_fetch_mmuBus_rsp_physicalAddress[25]
  PIN io_cpu_fetch_mmuBus_rsp_physicalAddress[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.630 246.000 482.910 250.000 ;
    END
  END io_cpu_fetch_mmuBus_rsp_physicalAddress[26]
  PIN io_cpu_fetch_mmuBus_rsp_physicalAddress[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.810 246.000 498.090 250.000 ;
    END
  END io_cpu_fetch_mmuBus_rsp_physicalAddress[27]
  PIN io_cpu_fetch_mmuBus_rsp_physicalAddress[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.990 246.000 513.270 250.000 ;
    END
  END io_cpu_fetch_mmuBus_rsp_physicalAddress[28]
  PIN io_cpu_fetch_mmuBus_rsp_physicalAddress[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 246.000 528.450 250.000 ;
    END
  END io_cpu_fetch_mmuBus_rsp_physicalAddress[29]
  PIN io_cpu_fetch_mmuBus_rsp_physicalAddress[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 246.000 104.790 250.000 ;
    END
  END io_cpu_fetch_mmuBus_rsp_physicalAddress[2]
  PIN io_cpu_fetch_mmuBus_rsp_physicalAddress[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.350 246.000 543.630 250.000 ;
    END
  END io_cpu_fetch_mmuBus_rsp_physicalAddress[30]
  PIN io_cpu_fetch_mmuBus_rsp_physicalAddress[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.530 246.000 558.810 250.000 ;
    END
  END io_cpu_fetch_mmuBus_rsp_physicalAddress[31]
  PIN io_cpu_fetch_mmuBus_rsp_physicalAddress[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.830 246.000 124.110 250.000 ;
    END
  END io_cpu_fetch_mmuBus_rsp_physicalAddress[3]
  PIN io_cpu_fetch_mmuBus_rsp_physicalAddress[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 246.000 140.670 250.000 ;
    END
  END io_cpu_fetch_mmuBus_rsp_physicalAddress[4]
  PIN io_cpu_fetch_mmuBus_rsp_physicalAddress[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 246.000 157.230 250.000 ;
    END
  END io_cpu_fetch_mmuBus_rsp_physicalAddress[5]
  PIN io_cpu_fetch_mmuBus_rsp_physicalAddress[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.510 246.000 173.790 250.000 ;
    END
  END io_cpu_fetch_mmuBus_rsp_physicalAddress[6]
  PIN io_cpu_fetch_mmuBus_rsp_physicalAddress[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 246.000 190.350 250.000 ;
    END
  END io_cpu_fetch_mmuBus_rsp_physicalAddress[7]
  PIN io_cpu_fetch_mmuBus_rsp_physicalAddress[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.630 246.000 206.910 250.000 ;
    END
  END io_cpu_fetch_mmuBus_rsp_physicalAddress[8]
  PIN io_cpu_fetch_mmuBus_rsp_physicalAddress[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 246.000 223.470 250.000 ;
    END
  END io_cpu_fetch_mmuBus_rsp_physicalAddress[9]
  PIN io_cpu_fetch_mmuBus_rsp_refilling
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 246.000 49.590 250.000 ;
    END
  END io_cpu_fetch_mmuBus_rsp_refilling
  PIN io_cpu_fetch_mmuBus_spr_payload_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 246.000 67.530 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_payload_data[0]
  PIN io_cpu_fetch_mmuBus_spr_payload_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.130 246.000 241.410 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_payload_data[10]
  PIN io_cpu_fetch_mmuBus_spr_payload_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.310 246.000 256.590 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_payload_data[11]
  PIN io_cpu_fetch_mmuBus_spr_payload_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.490 246.000 271.770 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_payload_data[12]
  PIN io_cpu_fetch_mmuBus_spr_payload_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 246.000 286.950 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_payload_data[13]
  PIN io_cpu_fetch_mmuBus_spr_payload_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 246.000 302.130 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_payload_data[14]
  PIN io_cpu_fetch_mmuBus_spr_payload_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.030 246.000 317.310 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_payload_data[15]
  PIN io_cpu_fetch_mmuBus_spr_payload_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.210 246.000 332.490 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_payload_data[16]
  PIN io_cpu_fetch_mmuBus_spr_payload_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 246.000 347.670 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_payload_data[17]
  PIN io_cpu_fetch_mmuBus_spr_payload_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.570 246.000 362.850 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_payload_data[18]
  PIN io_cpu_fetch_mmuBus_spr_payload_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.750 246.000 378.030 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_payload_data[19]
  PIN io_cpu_fetch_mmuBus_spr_payload_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 246.000 86.850 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_payload_data[1]
  PIN io_cpu_fetch_mmuBus_spr_payload_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 246.000 393.210 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_payload_data[20]
  PIN io_cpu_fetch_mmuBus_spr_payload_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.110 246.000 408.390 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_payload_data[21]
  PIN io_cpu_fetch_mmuBus_spr_payload_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.290 246.000 423.570 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_payload_data[22]
  PIN io_cpu_fetch_mmuBus_spr_payload_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.470 246.000 438.750 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_payload_data[23]
  PIN io_cpu_fetch_mmuBus_spr_payload_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.650 246.000 453.930 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_payload_data[24]
  PIN io_cpu_fetch_mmuBus_spr_payload_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.830 246.000 469.110 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_payload_data[25]
  PIN io_cpu_fetch_mmuBus_spr_payload_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.010 246.000 484.290 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_payload_data[26]
  PIN io_cpu_fetch_mmuBus_spr_payload_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 246.000 499.470 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_payload_data[27]
  PIN io_cpu_fetch_mmuBus_spr_payload_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.370 246.000 514.650 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_payload_data[28]
  PIN io_cpu_fetch_mmuBus_spr_payload_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.550 246.000 529.830 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_payload_data[29]
  PIN io_cpu_fetch_mmuBus_spr_payload_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 246.000 106.170 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_payload_data[2]
  PIN io_cpu_fetch_mmuBus_spr_payload_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.730 246.000 545.010 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_payload_data[30]
  PIN io_cpu_fetch_mmuBus_spr_payload_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.910 246.000 560.190 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_payload_data[31]
  PIN io_cpu_fetch_mmuBus_spr_payload_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.210 246.000 125.490 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_payload_data[3]
  PIN io_cpu_fetch_mmuBus_spr_payload_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 246.000 142.050 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_payload_data[4]
  PIN io_cpu_fetch_mmuBus_spr_payload_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.330 246.000 158.610 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_payload_data[5]
  PIN io_cpu_fetch_mmuBus_spr_payload_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 246.000 175.170 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_payload_data[6]
  PIN io_cpu_fetch_mmuBus_spr_payload_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 246.000 191.730 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_payload_data[7]
  PIN io_cpu_fetch_mmuBus_spr_payload_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.010 246.000 208.290 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_payload_data[8]
  PIN io_cpu_fetch_mmuBus_spr_payload_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 246.000 224.850 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_payload_data[9]
  PIN io_cpu_fetch_mmuBus_spr_payload_id[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 246.000 68.910 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_payload_id[0]
  PIN io_cpu_fetch_mmuBus_spr_payload_id[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 246.000 88.230 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_payload_id[1]
  PIN io_cpu_fetch_mmuBus_spr_payload_id[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 246.000 107.550 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_payload_id[2]
  PIN io_cpu_fetch_mmuBus_spr_payload_id[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 246.000 126.870 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_payload_id[3]
  PIN io_cpu_fetch_mmuBus_spr_payload_id[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.150 246.000 143.430 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_payload_id[4]
  PIN io_cpu_fetch_mmuBus_spr_payload_id[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.710 246.000 159.990 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_payload_id[5]
  PIN io_cpu_fetch_mmuBus_spr_payload_id[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 246.000 176.550 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_payload_id[6]
  PIN io_cpu_fetch_mmuBus_spr_payload_id[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.830 246.000 193.110 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_payload_id[7]
  PIN io_cpu_fetch_mmuBus_spr_payload_id[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 246.000 209.670 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_payload_id[8]
  PIN io_cpu_fetch_mmuBus_spr_payload_id[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.950 246.000 226.230 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_payload_id[9]
  PIN io_cpu_fetch_mmuBus_spr_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 246.000 50.970 250.000 ;
    END
  END io_cpu_fetch_mmuBus_spr_valid
  PIN io_cpu_fetch_pc[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 246.000 70.290 250.000 ;
    END
  END io_cpu_fetch_pc[0]
  PIN io_cpu_fetch_pc[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.510 246.000 242.790 250.000 ;
    END
  END io_cpu_fetch_pc[10]
  PIN io_cpu_fetch_pc[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 246.000 257.970 250.000 ;
    END
  END io_cpu_fetch_pc[11]
  PIN io_cpu_fetch_pc[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.870 246.000 273.150 250.000 ;
    END
  END io_cpu_fetch_pc[12]
  PIN io_cpu_fetch_pc[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 246.000 288.330 250.000 ;
    END
  END io_cpu_fetch_pc[13]
  PIN io_cpu_fetch_pc[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.230 246.000 303.510 250.000 ;
    END
  END io_cpu_fetch_pc[14]
  PIN io_cpu_fetch_pc[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.410 246.000 318.690 250.000 ;
    END
  END io_cpu_fetch_pc[15]
  PIN io_cpu_fetch_pc[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 246.000 333.870 250.000 ;
    END
  END io_cpu_fetch_pc[16]
  PIN io_cpu_fetch_pc[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.770 246.000 349.050 250.000 ;
    END
  END io_cpu_fetch_pc[17]
  PIN io_cpu_fetch_pc[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 246.000 364.230 250.000 ;
    END
  END io_cpu_fetch_pc[18]
  PIN io_cpu_fetch_pc[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.130 246.000 379.410 250.000 ;
    END
  END io_cpu_fetch_pc[19]
  PIN io_cpu_fetch_pc[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 246.000 89.610 250.000 ;
    END
  END io_cpu_fetch_pc[1]
  PIN io_cpu_fetch_pc[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.310 246.000 394.590 250.000 ;
    END
  END io_cpu_fetch_pc[20]
  PIN io_cpu_fetch_pc[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.490 246.000 409.770 250.000 ;
    END
  END io_cpu_fetch_pc[21]
  PIN io_cpu_fetch_pc[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.670 246.000 424.950 250.000 ;
    END
  END io_cpu_fetch_pc[22]
  PIN io_cpu_fetch_pc[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.850 246.000 440.130 250.000 ;
    END
  END io_cpu_fetch_pc[23]
  PIN io_cpu_fetch_pc[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.030 246.000 455.310 250.000 ;
    END
  END io_cpu_fetch_pc[24]
  PIN io_cpu_fetch_pc[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 246.000 470.490 250.000 ;
    END
  END io_cpu_fetch_pc[25]
  PIN io_cpu_fetch_pc[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.390 246.000 485.670 250.000 ;
    END
  END io_cpu_fetch_pc[26]
  PIN io_cpu_fetch_pc[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.570 246.000 500.850 250.000 ;
    END
  END io_cpu_fetch_pc[27]
  PIN io_cpu_fetch_pc[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.750 246.000 516.030 250.000 ;
    END
  END io_cpu_fetch_pc[28]
  PIN io_cpu_fetch_pc[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.930 246.000 531.210 250.000 ;
    END
  END io_cpu_fetch_pc[29]
  PIN io_cpu_fetch_pc[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 246.000 108.930 250.000 ;
    END
  END io_cpu_fetch_pc[2]
  PIN io_cpu_fetch_pc[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.110 246.000 546.390 250.000 ;
    END
  END io_cpu_fetch_pc[30]
  PIN io_cpu_fetch_pc[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.290 246.000 561.570 250.000 ;
    END
  END io_cpu_fetch_pc[31]
  PIN io_cpu_fetch_pc[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.970 246.000 128.250 250.000 ;
    END
  END io_cpu_fetch_pc[3]
  PIN io_cpu_fetch_pc[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 246.000 144.810 250.000 ;
    END
  END io_cpu_fetch_pc[4]
  PIN io_cpu_fetch_pc[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 246.000 161.370 250.000 ;
    END
  END io_cpu_fetch_pc[5]
  PIN io_cpu_fetch_pc[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 246.000 177.930 250.000 ;
    END
  END io_cpu_fetch_pc[6]
  PIN io_cpu_fetch_pc[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 246.000 194.490 250.000 ;
    END
  END io_cpu_fetch_pc[7]
  PIN io_cpu_fetch_pc[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.770 246.000 211.050 250.000 ;
    END
  END io_cpu_fetch_pc[8]
  PIN io_cpu_fetch_pc[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.330 246.000 227.610 250.000 ;
    END
  END io_cpu_fetch_pc[9]
  PIN io_cpu_fetch_physicalAddress[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 246.000 71.670 250.000 ;
    END
  END io_cpu_fetch_physicalAddress[0]
  PIN io_cpu_fetch_physicalAddress[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.890 246.000 244.170 250.000 ;
    END
  END io_cpu_fetch_physicalAddress[10]
  PIN io_cpu_fetch_physicalAddress[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.070 246.000 259.350 250.000 ;
    END
  END io_cpu_fetch_physicalAddress[11]
  PIN io_cpu_fetch_physicalAddress[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.250 246.000 274.530 250.000 ;
    END
  END io_cpu_fetch_physicalAddress[12]
  PIN io_cpu_fetch_physicalAddress[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.430 246.000 289.710 250.000 ;
    END
  END io_cpu_fetch_physicalAddress[13]
  PIN io_cpu_fetch_physicalAddress[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.610 246.000 304.890 250.000 ;
    END
  END io_cpu_fetch_physicalAddress[14]
  PIN io_cpu_fetch_physicalAddress[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 246.000 320.070 250.000 ;
    END
  END io_cpu_fetch_physicalAddress[15]
  PIN io_cpu_fetch_physicalAddress[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 246.000 335.250 250.000 ;
    END
  END io_cpu_fetch_physicalAddress[16]
  PIN io_cpu_fetch_physicalAddress[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.150 246.000 350.430 250.000 ;
    END
  END io_cpu_fetch_physicalAddress[17]
  PIN io_cpu_fetch_physicalAddress[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.330 246.000 365.610 250.000 ;
    END
  END io_cpu_fetch_physicalAddress[18]
  PIN io_cpu_fetch_physicalAddress[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.510 246.000 380.790 250.000 ;
    END
  END io_cpu_fetch_physicalAddress[19]
  PIN io_cpu_fetch_physicalAddress[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 246.000 90.990 250.000 ;
    END
  END io_cpu_fetch_physicalAddress[1]
  PIN io_cpu_fetch_physicalAddress[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.690 246.000 395.970 250.000 ;
    END
  END io_cpu_fetch_physicalAddress[20]
  PIN io_cpu_fetch_physicalAddress[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.870 246.000 411.150 250.000 ;
    END
  END io_cpu_fetch_physicalAddress[21]
  PIN io_cpu_fetch_physicalAddress[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.050 246.000 426.330 250.000 ;
    END
  END io_cpu_fetch_physicalAddress[22]
  PIN io_cpu_fetch_physicalAddress[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 246.000 441.510 250.000 ;
    END
  END io_cpu_fetch_physicalAddress[23]
  PIN io_cpu_fetch_physicalAddress[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.410 246.000 456.690 250.000 ;
    END
  END io_cpu_fetch_physicalAddress[24]
  PIN io_cpu_fetch_physicalAddress[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.590 246.000 471.870 250.000 ;
    END
  END io_cpu_fetch_physicalAddress[25]
  PIN io_cpu_fetch_physicalAddress[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.770 246.000 487.050 250.000 ;
    END
  END io_cpu_fetch_physicalAddress[26]
  PIN io_cpu_fetch_physicalAddress[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.950 246.000 502.230 250.000 ;
    END
  END io_cpu_fetch_physicalAddress[27]
  PIN io_cpu_fetch_physicalAddress[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.130 246.000 517.410 250.000 ;
    END
  END io_cpu_fetch_physicalAddress[28]
  PIN io_cpu_fetch_physicalAddress[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.310 246.000 532.590 250.000 ;
    END
  END io_cpu_fetch_physicalAddress[29]
  PIN io_cpu_fetch_physicalAddress[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 246.000 110.310 250.000 ;
    END
  END io_cpu_fetch_physicalAddress[2]
  PIN io_cpu_fetch_physicalAddress[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 246.000 547.770 250.000 ;
    END
  END io_cpu_fetch_physicalAddress[30]
  PIN io_cpu_fetch_physicalAddress[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.670 246.000 562.950 250.000 ;
    END
  END io_cpu_fetch_physicalAddress[31]
  PIN io_cpu_fetch_physicalAddress[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.350 246.000 129.630 250.000 ;
    END
  END io_cpu_fetch_physicalAddress[3]
  PIN io_cpu_fetch_physicalAddress[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 246.000 146.190 250.000 ;
    END
  END io_cpu_fetch_physicalAddress[4]
  PIN io_cpu_fetch_physicalAddress[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.470 246.000 162.750 250.000 ;
    END
  END io_cpu_fetch_physicalAddress[5]
  PIN io_cpu_fetch_physicalAddress[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.030 246.000 179.310 250.000 ;
    END
  END io_cpu_fetch_physicalAddress[6]
  PIN io_cpu_fetch_physicalAddress[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 246.000 195.870 250.000 ;
    END
  END io_cpu_fetch_physicalAddress[7]
  PIN io_cpu_fetch_physicalAddress[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.150 246.000 212.430 250.000 ;
    END
  END io_cpu_fetch_physicalAddress[8]
  PIN io_cpu_fetch_physicalAddress[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 246.000 228.990 250.000 ;
    END
  END io_cpu_fetch_physicalAddress[9]
  PIN io_cpu_fill_payload[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 246.000 73.050 250.000 ;
    END
  END io_cpu_fill_payload[0]
  PIN io_cpu_fill_payload[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.270 246.000 245.550 250.000 ;
    END
  END io_cpu_fill_payload[10]
  PIN io_cpu_fill_payload[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.450 246.000 260.730 250.000 ;
    END
  END io_cpu_fill_payload[11]
  PIN io_cpu_fill_payload[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.630 246.000 275.910 250.000 ;
    END
  END io_cpu_fill_payload[12]
  PIN io_cpu_fill_payload[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.810 246.000 291.090 250.000 ;
    END
  END io_cpu_fill_payload[13]
  PIN io_cpu_fill_payload[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 246.000 306.270 250.000 ;
    END
  END io_cpu_fill_payload[14]
  PIN io_cpu_fill_payload[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.170 246.000 321.450 250.000 ;
    END
  END io_cpu_fill_payload[15]
  PIN io_cpu_fill_payload[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.350 246.000 336.630 250.000 ;
    END
  END io_cpu_fill_payload[16]
  PIN io_cpu_fill_payload[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.530 246.000 351.810 250.000 ;
    END
  END io_cpu_fill_payload[17]
  PIN io_cpu_fill_payload[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.710 246.000 366.990 250.000 ;
    END
  END io_cpu_fill_payload[18]
  PIN io_cpu_fill_payload[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.890 246.000 382.170 250.000 ;
    END
  END io_cpu_fill_payload[19]
  PIN io_cpu_fill_payload[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 246.000 92.370 250.000 ;
    END
  END io_cpu_fill_payload[1]
  PIN io_cpu_fill_payload[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.070 246.000 397.350 250.000 ;
    END
  END io_cpu_fill_payload[20]
  PIN io_cpu_fill_payload[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 246.000 412.530 250.000 ;
    END
  END io_cpu_fill_payload[21]
  PIN io_cpu_fill_payload[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.430 246.000 427.710 250.000 ;
    END
  END io_cpu_fill_payload[22]
  PIN io_cpu_fill_payload[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.610 246.000 442.890 250.000 ;
    END
  END io_cpu_fill_payload[23]
  PIN io_cpu_fill_payload[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.790 246.000 458.070 250.000 ;
    END
  END io_cpu_fill_payload[24]
  PIN io_cpu_fill_payload[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.970 246.000 473.250 250.000 ;
    END
  END io_cpu_fill_payload[25]
  PIN io_cpu_fill_payload[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.150 246.000 488.430 250.000 ;
    END
  END io_cpu_fill_payload[26]
  PIN io_cpu_fill_payload[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.330 246.000 503.610 250.000 ;
    END
  END io_cpu_fill_payload[27]
  PIN io_cpu_fill_payload[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 246.000 518.790 250.000 ;
    END
  END io_cpu_fill_payload[28]
  PIN io_cpu_fill_payload[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.690 246.000 533.970 250.000 ;
    END
  END io_cpu_fill_payload[29]
  PIN io_cpu_fill_payload[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 246.000 111.690 250.000 ;
    END
  END io_cpu_fill_payload[2]
  PIN io_cpu_fill_payload[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.870 246.000 549.150 250.000 ;
    END
  END io_cpu_fill_payload[30]
  PIN io_cpu_fill_payload[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.050 246.000 564.330 250.000 ;
    END
  END io_cpu_fill_payload[31]
  PIN io_cpu_fill_payload[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.730 246.000 131.010 250.000 ;
    END
  END io_cpu_fill_payload[3]
  PIN io_cpu_fill_payload[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 246.000 147.570 250.000 ;
    END
  END io_cpu_fill_payload[4]
  PIN io_cpu_fill_payload[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.850 246.000 164.130 250.000 ;
    END
  END io_cpu_fill_payload[5]
  PIN io_cpu_fill_payload[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 246.000 180.690 250.000 ;
    END
  END io_cpu_fill_payload[6]
  PIN io_cpu_fill_payload[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 246.000 197.250 250.000 ;
    END
  END io_cpu_fill_payload[7]
  PIN io_cpu_fill_payload[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.530 246.000 213.810 250.000 ;
    END
  END io_cpu_fill_payload[8]
  PIN io_cpu_fill_payload[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.090 246.000 230.370 250.000 ;
    END
  END io_cpu_fill_payload[9]
  PIN io_cpu_fill_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 246.000 52.350 250.000 ;
    END
  END io_cpu_fill_valid
  PIN io_cpu_prefetch_haltIt
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 246.000 53.730 250.000 ;
    END
  END io_cpu_prefetch_haltIt
  PIN io_cpu_prefetch_isValid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 246.000 55.110 250.000 ;
    END
  END io_cpu_prefetch_isValid
  PIN io_cpu_prefetch_pc[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 246.000 74.430 250.000 ;
    END
  END io_cpu_prefetch_pc[0]
  PIN io_cpu_prefetch_pc[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 246.000 246.930 250.000 ;
    END
  END io_cpu_prefetch_pc[10]
  PIN io_cpu_prefetch_pc[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 246.000 262.110 250.000 ;
    END
  END io_cpu_prefetch_pc[11]
  PIN io_cpu_prefetch_pc[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 246.000 277.290 250.000 ;
    END
  END io_cpu_prefetch_pc[12]
  PIN io_cpu_prefetch_pc[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 246.000 292.470 250.000 ;
    END
  END io_cpu_prefetch_pc[13]
  PIN io_cpu_prefetch_pc[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.370 246.000 307.650 250.000 ;
    END
  END io_cpu_prefetch_pc[14]
  PIN io_cpu_prefetch_pc[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 246.000 322.830 250.000 ;
    END
  END io_cpu_prefetch_pc[15]
  PIN io_cpu_prefetch_pc[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.730 246.000 338.010 250.000 ;
    END
  END io_cpu_prefetch_pc[16]
  PIN io_cpu_prefetch_pc[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.910 246.000 353.190 250.000 ;
    END
  END io_cpu_prefetch_pc[17]
  PIN io_cpu_prefetch_pc[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.090 246.000 368.370 250.000 ;
    END
  END io_cpu_prefetch_pc[18]
  PIN io_cpu_prefetch_pc[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 246.000 383.550 250.000 ;
    END
  END io_cpu_prefetch_pc[19]
  PIN io_cpu_prefetch_pc[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 246.000 93.750 250.000 ;
    END
  END io_cpu_prefetch_pc[1]
  PIN io_cpu_prefetch_pc[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.450 246.000 398.730 250.000 ;
    END
  END io_cpu_prefetch_pc[20]
  PIN io_cpu_prefetch_pc[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.630 246.000 413.910 250.000 ;
    END
  END io_cpu_prefetch_pc[21]
  PIN io_cpu_prefetch_pc[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.810 246.000 429.090 250.000 ;
    END
  END io_cpu_prefetch_pc[22]
  PIN io_cpu_prefetch_pc[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.990 246.000 444.270 250.000 ;
    END
  END io_cpu_prefetch_pc[23]
  PIN io_cpu_prefetch_pc[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.170 246.000 459.450 250.000 ;
    END
  END io_cpu_prefetch_pc[24]
  PIN io_cpu_prefetch_pc[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.350 246.000 474.630 250.000 ;
    END
  END io_cpu_prefetch_pc[25]
  PIN io_cpu_prefetch_pc[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 246.000 489.810 250.000 ;
    END
  END io_cpu_prefetch_pc[26]
  PIN io_cpu_prefetch_pc[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.710 246.000 504.990 250.000 ;
    END
  END io_cpu_prefetch_pc[27]
  PIN io_cpu_prefetch_pc[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.890 246.000 520.170 250.000 ;
    END
  END io_cpu_prefetch_pc[28]
  PIN io_cpu_prefetch_pc[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.070 246.000 535.350 250.000 ;
    END
  END io_cpu_prefetch_pc[29]
  PIN io_cpu_prefetch_pc[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 246.000 113.070 250.000 ;
    END
  END io_cpu_prefetch_pc[2]
  PIN io_cpu_prefetch_pc[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.250 246.000 550.530 250.000 ;
    END
  END io_cpu_prefetch_pc[30]
  PIN io_cpu_prefetch_pc[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.430 246.000 565.710 250.000 ;
    END
  END io_cpu_prefetch_pc[31]
  PIN io_cpu_prefetch_pc[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 246.000 132.390 250.000 ;
    END
  END io_cpu_prefetch_pc[3]
  PIN io_cpu_prefetch_pc[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.670 246.000 148.950 250.000 ;
    END
  END io_cpu_prefetch_pc[4]
  PIN io_cpu_prefetch_pc[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.230 246.000 165.510 250.000 ;
    END
  END io_cpu_prefetch_pc[5]
  PIN io_cpu_prefetch_pc[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 246.000 182.070 250.000 ;
    END
  END io_cpu_prefetch_pc[6]
  PIN io_cpu_prefetch_pc[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.350 246.000 198.630 250.000 ;
    END
  END io_cpu_prefetch_pc[7]
  PIN io_cpu_prefetch_pc[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 246.000 215.190 250.000 ;
    END
  END io_cpu_prefetch_pc[8]
  PIN io_cpu_prefetch_pc[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.470 246.000 231.750 250.000 ;
    END
  END io_cpu_prefetch_pc[9]
  PIN io_flush
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 246.000 567.090 250.000 ;
    END
  END io_flush
  PIN io_mem_cmd_payload_address[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 4.000 ;
    END
  END io_mem_cmd_payload_address[0]
  PIN io_mem_cmd_payload_address[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 0.000 255.210 4.000 ;
    END
  END io_mem_cmd_payload_address[10]
  PIN io_mem_cmd_payload_address[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.410 0.000 272.690 4.000 ;
    END
  END io_mem_cmd_payload_address[11]
  PIN io_mem_cmd_payload_address[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END io_mem_cmd_payload_address[12]
  PIN io_mem_cmd_payload_address[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.370 0.000 307.650 4.000 ;
    END
  END io_mem_cmd_payload_address[13]
  PIN io_mem_cmd_payload_address[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.850 0.000 325.130 4.000 ;
    END
  END io_mem_cmd_payload_address[14]
  PIN io_mem_cmd_payload_address[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.330 0.000 342.610 4.000 ;
    END
  END io_mem_cmd_payload_address[15]
  PIN io_mem_cmd_payload_address[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.810 0.000 360.090 4.000 ;
    END
  END io_mem_cmd_payload_address[16]
  PIN io_mem_cmd_payload_address[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 0.000 377.570 4.000 ;
    END
  END io_mem_cmd_payload_address[17]
  PIN io_mem_cmd_payload_address[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.770 0.000 395.050 4.000 ;
    END
  END io_mem_cmd_payload_address[18]
  PIN io_mem_cmd_payload_address[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END io_mem_cmd_payload_address[19]
  PIN io_mem_cmd_payload_address[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 4.000 ;
    END
  END io_mem_cmd_payload_address[1]
  PIN io_mem_cmd_payload_address[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.730 0.000 430.010 4.000 ;
    END
  END io_mem_cmd_payload_address[20]
  PIN io_mem_cmd_payload_address[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.210 0.000 447.490 4.000 ;
    END
  END io_mem_cmd_payload_address[21]
  PIN io_mem_cmd_payload_address[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.690 0.000 464.970 4.000 ;
    END
  END io_mem_cmd_payload_address[22]
  PIN io_mem_cmd_payload_address[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.170 0.000 482.450 4.000 ;
    END
  END io_mem_cmd_payload_address[23]
  PIN io_mem_cmd_payload_address[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.650 0.000 499.930 4.000 ;
    END
  END io_mem_cmd_payload_address[24]
  PIN io_mem_cmd_payload_address[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.130 0.000 517.410 4.000 ;
    END
  END io_mem_cmd_payload_address[25]
  PIN io_mem_cmd_payload_address[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 0.000 534.890 4.000 ;
    END
  END io_mem_cmd_payload_address[26]
  PIN io_mem_cmd_payload_address[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.090 0.000 552.370 4.000 ;
    END
  END io_mem_cmd_payload_address[27]
  PIN io_mem_cmd_payload_address[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.570 0.000 569.850 4.000 ;
    END
  END io_mem_cmd_payload_address[28]
  PIN io_mem_cmd_payload_address[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.050 0.000 587.330 4.000 ;
    END
  END io_mem_cmd_payload_address[29]
  PIN io_mem_cmd_payload_address[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END io_mem_cmd_payload_address[2]
  PIN io_mem_cmd_payload_address[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.530 0.000 604.810 4.000 ;
    END
  END io_mem_cmd_payload_address[30]
  PIN io_mem_cmd_payload_address[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.010 0.000 622.290 4.000 ;
    END
  END io_mem_cmd_payload_address[31]
  PIN io_mem_cmd_payload_address[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 4.000 ;
    END
  END io_mem_cmd_payload_address[3]
  PIN io_mem_cmd_payload_address[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 4.000 ;
    END
  END io_mem_cmd_payload_address[4]
  PIN io_mem_cmd_payload_address[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END io_mem_cmd_payload_address[5]
  PIN io_mem_cmd_payload_address[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 4.000 ;
    END
  END io_mem_cmd_payload_address[6]
  PIN io_mem_cmd_payload_address[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.490 0.000 202.770 4.000 ;
    END
  END io_mem_cmd_payload_address[7]
  PIN io_mem_cmd_payload_address[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.970 0.000 220.250 4.000 ;
    END
  END io_mem_cmd_payload_address[8]
  PIN io_mem_cmd_payload_address[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 0.000 237.730 4.000 ;
    END
  END io_mem_cmd_payload_address[9]
  PIN io_mem_cmd_payload_size[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END io_mem_cmd_payload_size[0]
  PIN io_mem_cmd_payload_size[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 0.000 89.150 4.000 ;
    END
  END io_mem_cmd_payload_size[1]
  PIN io_mem_cmd_payload_size[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END io_mem_cmd_payload_size[2]
  PIN io_mem_cmd_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 0.000 19.230 4.000 ;
    END
  END io_mem_cmd_ready
  PIN io_mem_cmd_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END io_mem_cmd_valid
  PIN io_mem_rsp_payload_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 4.000 ;
    END
  END io_mem_rsp_payload_data[0]
  PIN io_mem_rsp_payload_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 0.000 263.950 4.000 ;
    END
  END io_mem_rsp_payload_data[10]
  PIN io_mem_rsp_payload_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 0.000 281.430 4.000 ;
    END
  END io_mem_rsp_payload_data[11]
  PIN io_mem_rsp_payload_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.630 0.000 298.910 4.000 ;
    END
  END io_mem_rsp_payload_data[12]
  PIN io_mem_rsp_payload_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.110 0.000 316.390 4.000 ;
    END
  END io_mem_rsp_payload_data[13]
  PIN io_mem_rsp_payload_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 0.000 333.870 4.000 ;
    END
  END io_mem_rsp_payload_data[14]
  PIN io_mem_rsp_payload_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 4.000 ;
    END
  END io_mem_rsp_payload_data[15]
  PIN io_mem_rsp_payload_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.550 0.000 368.830 4.000 ;
    END
  END io_mem_rsp_payload_data[16]
  PIN io_mem_rsp_payload_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.030 0.000 386.310 4.000 ;
    END
  END io_mem_rsp_payload_data[17]
  PIN io_mem_rsp_payload_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.510 0.000 403.790 4.000 ;
    END
  END io_mem_rsp_payload_data[18]
  PIN io_mem_rsp_payload_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.990 0.000 421.270 4.000 ;
    END
  END io_mem_rsp_payload_data[19]
  PIN io_mem_rsp_payload_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 4.000 ;
    END
  END io_mem_rsp_payload_data[1]
  PIN io_mem_rsp_payload_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.470 0.000 438.750 4.000 ;
    END
  END io_mem_rsp_payload_data[20]
  PIN io_mem_rsp_payload_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.950 0.000 456.230 4.000 ;
    END
  END io_mem_rsp_payload_data[21]
  PIN io_mem_rsp_payload_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 0.000 473.710 4.000 ;
    END
  END io_mem_rsp_payload_data[22]
  PIN io_mem_rsp_payload_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.910 0.000 491.190 4.000 ;
    END
  END io_mem_rsp_payload_data[23]
  PIN io_mem_rsp_payload_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.390 0.000 508.670 4.000 ;
    END
  END io_mem_rsp_payload_data[24]
  PIN io_mem_rsp_payload_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.870 0.000 526.150 4.000 ;
    END
  END io_mem_rsp_payload_data[25]
  PIN io_mem_rsp_payload_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.350 0.000 543.630 4.000 ;
    END
  END io_mem_rsp_payload_data[26]
  PIN io_mem_rsp_payload_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.830 0.000 561.110 4.000 ;
    END
  END io_mem_rsp_payload_data[27]
  PIN io_mem_rsp_payload_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.310 0.000 578.590 4.000 ;
    END
  END io_mem_rsp_payload_data[28]
  PIN io_mem_rsp_payload_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 0.000 596.070 4.000 ;
    END
  END io_mem_rsp_payload_data[29]
  PIN io_mem_rsp_payload_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.830 0.000 124.110 4.000 ;
    END
  END io_mem_rsp_payload_data[2]
  PIN io_mem_rsp_payload_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.270 0.000 613.550 4.000 ;
    END
  END io_mem_rsp_payload_data[30]
  PIN io_mem_rsp_payload_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.750 0.000 631.030 4.000 ;
    END
  END io_mem_rsp_payload_data[31]
  PIN io_mem_rsp_payload_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.310 0.000 141.590 4.000 ;
    END
  END io_mem_rsp_payload_data[3]
  PIN io_mem_rsp_payload_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 0.000 159.070 4.000 ;
    END
  END io_mem_rsp_payload_data[4]
  PIN io_mem_rsp_payload_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 0.000 176.550 4.000 ;
    END
  END io_mem_rsp_payload_data[5]
  PIN io_mem_rsp_payload_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.750 0.000 194.030 4.000 ;
    END
  END io_mem_rsp_payload_data[6]
  PIN io_mem_rsp_payload_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 0.000 211.510 4.000 ;
    END
  END io_mem_rsp_payload_data[7]
  PIN io_mem_rsp_payload_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END io_mem_rsp_payload_data[8]
  PIN io_mem_rsp_payload_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.190 0.000 246.470 4.000 ;
    END
  END io_mem_rsp_payload_data[9]
  PIN io_mem_rsp_payload_error
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 4.000 ;
    END
  END io_mem_rsp_payload_error
  PIN io_mem_rsp_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END io_mem_rsp_valid
  PIN io_spr_payload_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.570 246.000 569.850 250.000 ;
    END
  END io_spr_payload_data[0]
  PIN io_spr_payload_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.170 246.000 597.450 250.000 ;
    END
  END io_spr_payload_data[10]
  PIN io_spr_payload_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.550 246.000 598.830 250.000 ;
    END
  END io_spr_payload_data[11]
  PIN io_spr_payload_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.930 246.000 600.210 250.000 ;
    END
  END io_spr_payload_data[12]
  PIN io_spr_payload_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.310 246.000 601.590 250.000 ;
    END
  END io_spr_payload_data[13]
  PIN io_spr_payload_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.690 246.000 602.970 250.000 ;
    END
  END io_spr_payload_data[14]
  PIN io_spr_payload_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.070 246.000 604.350 250.000 ;
    END
  END io_spr_payload_data[15]
  PIN io_spr_payload_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.450 246.000 605.730 250.000 ;
    END
  END io_spr_payload_data[16]
  PIN io_spr_payload_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.830 246.000 607.110 250.000 ;
    END
  END io_spr_payload_data[17]
  PIN io_spr_payload_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.210 246.000 608.490 250.000 ;
    END
  END io_spr_payload_data[18]
  PIN io_spr_payload_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.590 246.000 609.870 250.000 ;
    END
  END io_spr_payload_data[19]
  PIN io_spr_payload_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.330 246.000 572.610 250.000 ;
    END
  END io_spr_payload_data[1]
  PIN io_spr_payload_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.970 246.000 611.250 250.000 ;
    END
  END io_spr_payload_data[20]
  PIN io_spr_payload_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.350 246.000 612.630 250.000 ;
    END
  END io_spr_payload_data[21]
  PIN io_spr_payload_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.730 246.000 614.010 250.000 ;
    END
  END io_spr_payload_data[22]
  PIN io_spr_payload_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.110 246.000 615.390 250.000 ;
    END
  END io_spr_payload_data[23]
  PIN io_spr_payload_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.490 246.000 616.770 250.000 ;
    END
  END io_spr_payload_data[24]
  PIN io_spr_payload_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.870 246.000 618.150 250.000 ;
    END
  END io_spr_payload_data[25]
  PIN io_spr_payload_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.250 246.000 619.530 250.000 ;
    END
  END io_spr_payload_data[26]
  PIN io_spr_payload_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.630 246.000 620.910 250.000 ;
    END
  END io_spr_payload_data[27]
  PIN io_spr_payload_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.010 246.000 622.290 250.000 ;
    END
  END io_spr_payload_data[28]
  PIN io_spr_payload_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.390 246.000 623.670 250.000 ;
    END
  END io_spr_payload_data[29]
  PIN io_spr_payload_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.090 246.000 575.370 250.000 ;
    END
  END io_spr_payload_data[2]
  PIN io_spr_payload_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 246.000 625.050 250.000 ;
    END
  END io_spr_payload_data[30]
  PIN io_spr_payload_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.150 246.000 626.430 250.000 ;
    END
  END io_spr_payload_data[31]
  PIN io_spr_payload_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.850 246.000 578.130 250.000 ;
    END
  END io_spr_payload_data[3]
  PIN io_spr_payload_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.610 246.000 580.890 250.000 ;
    END
  END io_spr_payload_data[4]
  PIN io_spr_payload_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.370 246.000 583.650 250.000 ;
    END
  END io_spr_payload_data[5]
  PIN io_spr_payload_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.130 246.000 586.410 250.000 ;
    END
  END io_spr_payload_data[6]
  PIN io_spr_payload_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.890 246.000 589.170 250.000 ;
    END
  END io_spr_payload_data[7]
  PIN io_spr_payload_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.650 246.000 591.930 250.000 ;
    END
  END io_spr_payload_data[8]
  PIN io_spr_payload_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.410 246.000 594.690 250.000 ;
    END
  END io_spr_payload_data[9]
  PIN io_spr_payload_id[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.950 246.000 571.230 250.000 ;
    END
  END io_spr_payload_id[0]
  PIN io_spr_payload_id[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.710 246.000 573.990 250.000 ;
    END
  END io_spr_payload_id[1]
  PIN io_spr_payload_id[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.470 246.000 576.750 250.000 ;
    END
  END io_spr_payload_id[2]
  PIN io_spr_payload_id[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.230 246.000 579.510 250.000 ;
    END
  END io_spr_payload_id[3]
  PIN io_spr_payload_id[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.990 246.000 582.270 250.000 ;
    END
  END io_spr_payload_id[4]
  PIN io_spr_payload_id[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.750 246.000 585.030 250.000 ;
    END
  END io_spr_payload_id[5]
  PIN io_spr_payload_id[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.510 246.000 587.790 250.000 ;
    END
  END io_spr_payload_id[6]
  PIN io_spr_payload_id[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.270 246.000 590.550 250.000 ;
    END
  END io_spr_payload_id[7]
  PIN io_spr_payload_id[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.030 246.000 593.310 250.000 ;
    END
  END io_spr_payload_id[8]
  PIN io_spr_payload_id[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 246.000 596.070 250.000 ;
    END
  END io_spr_payload_id[9]
  PIN io_spr_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.190 246.000 568.470 250.000 ;
    END
  END io_spr_valid
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.910 246.000 629.190 250.000 ;
    END
  END reset
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 179.160 22.640 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 179.160 176.240 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 179.160 329.840 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 179.160 483.440 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 7.940 10.640 9.540 182.480 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 179.160 99.440 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 179.160 253.040 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 179.160 406.640 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 179.160 560.240 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 10.700 10.640 12.300 182.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 630.780 10.640 632.380 179.760 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 235.225 644.650 236.830 ;
        RECT 5.330 229.785 644.650 232.615 ;
        RECT 5.330 224.345 644.650 227.175 ;
        RECT 5.330 218.905 644.650 221.735 ;
        RECT 5.330 213.465 644.650 216.295 ;
        RECT 5.330 208.025 644.650 210.855 ;
        RECT 5.330 202.585 644.650 205.415 ;
        RECT 5.330 197.145 644.650 199.975 ;
        RECT 5.330 191.705 644.650 194.535 ;
        RECT 5.330 186.265 644.650 189.095 ;
        RECT 5.330 180.825 644.650 183.655 ;
        RECT 5.330 175.385 14.910 178.215 ;
        RECT 5.330 169.945 14.910 172.775 ;
        RECT 5.330 164.505 14.910 167.335 ;
        RECT 5.330 159.065 14.910 161.895 ;
        RECT 5.330 153.625 14.910 156.455 ;
        RECT 5.330 148.185 14.910 151.015 ;
        RECT 5.330 142.745 14.910 145.575 ;
        RECT 5.330 137.305 14.910 140.135 ;
        RECT 5.330 131.865 14.910 134.695 ;
        RECT 5.330 126.425 14.910 129.255 ;
        RECT 5.330 120.985 14.910 123.815 ;
        RECT 5.330 115.545 14.910 118.375 ;
        RECT 5.330 110.105 14.910 112.935 ;
        RECT 5.330 104.665 14.910 107.495 ;
        RECT 5.330 99.225 14.910 102.055 ;
        RECT 5.330 93.785 14.910 96.615 ;
        RECT 5.330 88.345 14.910 91.175 ;
        RECT 5.330 82.905 14.910 85.735 ;
        RECT 5.330 77.465 14.910 80.295 ;
        RECT 5.330 72.025 14.910 74.855 ;
        RECT 5.330 66.585 14.910 69.415 ;
        RECT 5.330 61.145 14.910 63.975 ;
        RECT 5.330 55.705 14.910 58.535 ;
        RECT 5.330 50.265 14.910 53.095 ;
        RECT 5.330 44.825 14.910 47.655 ;
        RECT 5.330 39.385 14.910 42.215 ;
        RECT 5.330 33.945 14.910 36.775 ;
        RECT 5.330 28.505 14.910 31.335 ;
        RECT 5.330 23.065 14.910 25.895 ;
        RECT 5.330 17.625 14.910 20.455 ;
        RECT 5.330 13.790 14.910 15.015 ;
        RECT 5.330 12.185 644.650 13.790 ;
      LAYER li1 ;
        RECT 5.520 10.795 644.460 236.725 ;
      LAYER met1 ;
        RECT 5.520 9.220 644.460 249.860 ;
      LAYER met2 ;
        RECT 7.970 245.720 20.050 249.970 ;
        RECT 20.890 245.720 21.430 249.970 ;
        RECT 22.270 245.720 22.810 249.970 ;
        RECT 23.650 245.720 24.190 249.970 ;
        RECT 25.030 245.720 25.570 249.970 ;
        RECT 26.410 245.720 26.950 249.970 ;
        RECT 27.790 245.720 28.330 249.970 ;
        RECT 29.170 245.720 29.710 249.970 ;
        RECT 30.550 245.720 31.090 249.970 ;
        RECT 31.930 245.720 32.470 249.970 ;
        RECT 33.310 245.720 33.850 249.970 ;
        RECT 34.690 245.720 35.230 249.970 ;
        RECT 36.070 245.720 36.610 249.970 ;
        RECT 37.450 245.720 37.990 249.970 ;
        RECT 38.830 245.720 39.370 249.970 ;
        RECT 40.210 245.720 40.750 249.970 ;
        RECT 41.590 245.720 42.130 249.970 ;
        RECT 42.970 245.720 43.510 249.970 ;
        RECT 44.350 245.720 44.890 249.970 ;
        RECT 45.730 245.720 46.270 249.970 ;
        RECT 47.110 245.720 47.650 249.970 ;
        RECT 48.490 245.720 49.030 249.970 ;
        RECT 49.870 245.720 50.410 249.970 ;
        RECT 51.250 245.720 51.790 249.970 ;
        RECT 52.630 245.720 53.170 249.970 ;
        RECT 54.010 245.720 54.550 249.970 ;
        RECT 55.390 245.720 55.930 249.970 ;
        RECT 56.770 245.720 57.310 249.970 ;
        RECT 58.150 245.720 58.690 249.970 ;
        RECT 59.530 245.720 60.070 249.970 ;
        RECT 60.910 245.720 61.450 249.970 ;
        RECT 62.290 245.720 62.830 249.970 ;
        RECT 63.670 245.720 64.210 249.970 ;
        RECT 65.050 245.720 65.590 249.970 ;
        RECT 66.430 245.720 66.970 249.970 ;
        RECT 67.810 245.720 68.350 249.970 ;
        RECT 69.190 245.720 69.730 249.970 ;
        RECT 70.570 245.720 71.110 249.970 ;
        RECT 71.950 245.720 72.490 249.970 ;
        RECT 73.330 245.720 73.870 249.970 ;
        RECT 74.710 245.720 75.250 249.970 ;
        RECT 76.090 245.720 76.630 249.970 ;
        RECT 77.470 245.720 78.010 249.970 ;
        RECT 78.850 245.720 79.390 249.970 ;
        RECT 80.230 245.720 80.770 249.970 ;
        RECT 81.610 245.720 82.150 249.970 ;
        RECT 82.990 245.720 83.530 249.970 ;
        RECT 84.370 245.720 84.910 249.970 ;
        RECT 85.750 245.720 86.290 249.970 ;
        RECT 87.130 245.720 87.670 249.970 ;
        RECT 88.510 245.720 89.050 249.970 ;
        RECT 89.890 245.720 90.430 249.970 ;
        RECT 91.270 245.720 91.810 249.970 ;
        RECT 92.650 245.720 93.190 249.970 ;
        RECT 94.030 245.720 94.570 249.970 ;
        RECT 95.410 245.720 95.950 249.970 ;
        RECT 96.790 245.720 97.330 249.970 ;
        RECT 98.170 245.720 98.710 249.970 ;
        RECT 99.550 245.720 100.090 249.970 ;
        RECT 100.930 245.720 101.470 249.970 ;
        RECT 102.310 245.720 102.850 249.970 ;
        RECT 103.690 245.720 104.230 249.970 ;
        RECT 105.070 245.720 105.610 249.970 ;
        RECT 106.450 245.720 106.990 249.970 ;
        RECT 107.830 245.720 108.370 249.970 ;
        RECT 109.210 245.720 109.750 249.970 ;
        RECT 110.590 245.720 111.130 249.970 ;
        RECT 111.970 245.720 112.510 249.970 ;
        RECT 113.350 245.720 113.890 249.970 ;
        RECT 114.730 245.720 115.270 249.970 ;
        RECT 116.110 245.720 116.650 249.970 ;
        RECT 117.490 245.720 118.030 249.970 ;
        RECT 118.870 245.720 119.410 249.970 ;
        RECT 120.250 245.720 120.790 249.970 ;
        RECT 121.630 245.720 122.170 249.970 ;
        RECT 123.010 245.720 123.550 249.970 ;
        RECT 124.390 245.720 124.930 249.970 ;
        RECT 125.770 245.720 126.310 249.970 ;
        RECT 127.150 245.720 127.690 249.970 ;
        RECT 128.530 245.720 129.070 249.970 ;
        RECT 129.910 245.720 130.450 249.970 ;
        RECT 131.290 245.720 131.830 249.970 ;
        RECT 132.670 245.720 133.210 249.970 ;
        RECT 134.050 245.720 134.590 249.970 ;
        RECT 135.430 245.720 135.970 249.970 ;
        RECT 136.810 245.720 137.350 249.970 ;
        RECT 138.190 245.720 138.730 249.970 ;
        RECT 139.570 245.720 140.110 249.970 ;
        RECT 140.950 245.720 141.490 249.970 ;
        RECT 142.330 245.720 142.870 249.970 ;
        RECT 143.710 245.720 144.250 249.970 ;
        RECT 145.090 245.720 145.630 249.970 ;
        RECT 146.470 245.720 147.010 249.970 ;
        RECT 147.850 245.720 148.390 249.970 ;
        RECT 149.230 245.720 149.770 249.970 ;
        RECT 150.610 245.720 151.150 249.970 ;
        RECT 151.990 245.720 152.530 249.970 ;
        RECT 153.370 245.720 153.910 249.970 ;
        RECT 154.750 245.720 155.290 249.970 ;
        RECT 156.130 245.720 156.670 249.970 ;
        RECT 157.510 245.720 158.050 249.970 ;
        RECT 158.890 245.720 159.430 249.970 ;
        RECT 160.270 245.720 160.810 249.970 ;
        RECT 161.650 245.720 162.190 249.970 ;
        RECT 163.030 245.720 163.570 249.970 ;
        RECT 164.410 245.720 164.950 249.970 ;
        RECT 165.790 245.720 166.330 249.970 ;
        RECT 167.170 245.720 167.710 249.970 ;
        RECT 168.550 245.720 169.090 249.970 ;
        RECT 169.930 245.720 170.470 249.970 ;
        RECT 171.310 245.720 171.850 249.970 ;
        RECT 172.690 245.720 173.230 249.970 ;
        RECT 174.070 245.720 174.610 249.970 ;
        RECT 175.450 245.720 175.990 249.970 ;
        RECT 176.830 245.720 177.370 249.970 ;
        RECT 178.210 245.720 178.750 249.970 ;
        RECT 179.590 245.720 180.130 249.970 ;
        RECT 180.970 245.720 181.510 249.970 ;
        RECT 182.350 245.720 182.890 249.970 ;
        RECT 183.730 245.720 184.270 249.970 ;
        RECT 185.110 245.720 185.650 249.970 ;
        RECT 186.490 245.720 187.030 249.970 ;
        RECT 187.870 245.720 188.410 249.970 ;
        RECT 189.250 245.720 189.790 249.970 ;
        RECT 190.630 245.720 191.170 249.970 ;
        RECT 192.010 245.720 192.550 249.970 ;
        RECT 193.390 245.720 193.930 249.970 ;
        RECT 194.770 245.720 195.310 249.970 ;
        RECT 196.150 245.720 196.690 249.970 ;
        RECT 197.530 245.720 198.070 249.970 ;
        RECT 198.910 245.720 199.450 249.970 ;
        RECT 200.290 245.720 200.830 249.970 ;
        RECT 201.670 245.720 202.210 249.970 ;
        RECT 203.050 245.720 203.590 249.970 ;
        RECT 204.430 245.720 204.970 249.970 ;
        RECT 205.810 245.720 206.350 249.970 ;
        RECT 207.190 245.720 207.730 249.970 ;
        RECT 208.570 245.720 209.110 249.970 ;
        RECT 209.950 245.720 210.490 249.970 ;
        RECT 211.330 245.720 211.870 249.970 ;
        RECT 212.710 245.720 213.250 249.970 ;
        RECT 214.090 245.720 214.630 249.970 ;
        RECT 215.470 245.720 216.010 249.970 ;
        RECT 216.850 245.720 217.390 249.970 ;
        RECT 218.230 245.720 218.770 249.970 ;
        RECT 219.610 245.720 220.150 249.970 ;
        RECT 220.990 245.720 221.530 249.970 ;
        RECT 222.370 245.720 222.910 249.970 ;
        RECT 223.750 245.720 224.290 249.970 ;
        RECT 225.130 245.720 225.670 249.970 ;
        RECT 226.510 245.720 227.050 249.970 ;
        RECT 227.890 245.720 228.430 249.970 ;
        RECT 229.270 245.720 229.810 249.970 ;
        RECT 230.650 245.720 231.190 249.970 ;
        RECT 232.030 245.720 232.570 249.970 ;
        RECT 233.410 245.720 233.950 249.970 ;
        RECT 234.790 245.720 235.330 249.970 ;
        RECT 236.170 245.720 236.710 249.970 ;
        RECT 237.550 245.720 238.090 249.970 ;
        RECT 238.930 245.720 239.470 249.970 ;
        RECT 240.310 245.720 240.850 249.970 ;
        RECT 241.690 245.720 242.230 249.970 ;
        RECT 243.070 245.720 243.610 249.970 ;
        RECT 244.450 245.720 244.990 249.970 ;
        RECT 245.830 245.720 246.370 249.970 ;
        RECT 247.210 245.720 247.750 249.970 ;
        RECT 248.590 245.720 249.130 249.970 ;
        RECT 249.970 245.720 250.510 249.970 ;
        RECT 251.350 245.720 251.890 249.970 ;
        RECT 252.730 245.720 253.270 249.970 ;
        RECT 254.110 245.720 254.650 249.970 ;
        RECT 255.490 245.720 256.030 249.970 ;
        RECT 256.870 245.720 257.410 249.970 ;
        RECT 258.250 245.720 258.790 249.970 ;
        RECT 259.630 245.720 260.170 249.970 ;
        RECT 261.010 245.720 261.550 249.970 ;
        RECT 262.390 245.720 262.930 249.970 ;
        RECT 263.770 245.720 264.310 249.970 ;
        RECT 265.150 245.720 265.690 249.970 ;
        RECT 266.530 245.720 267.070 249.970 ;
        RECT 267.910 245.720 268.450 249.970 ;
        RECT 269.290 245.720 269.830 249.970 ;
        RECT 270.670 245.720 271.210 249.970 ;
        RECT 272.050 245.720 272.590 249.970 ;
        RECT 273.430 245.720 273.970 249.970 ;
        RECT 274.810 245.720 275.350 249.970 ;
        RECT 276.190 245.720 276.730 249.970 ;
        RECT 277.570 245.720 278.110 249.970 ;
        RECT 278.950 245.720 279.490 249.970 ;
        RECT 280.330 245.720 280.870 249.970 ;
        RECT 281.710 245.720 282.250 249.970 ;
        RECT 283.090 245.720 283.630 249.970 ;
        RECT 284.470 245.720 285.010 249.970 ;
        RECT 285.850 245.720 286.390 249.970 ;
        RECT 287.230 245.720 287.770 249.970 ;
        RECT 288.610 245.720 289.150 249.970 ;
        RECT 289.990 245.720 290.530 249.970 ;
        RECT 291.370 245.720 291.910 249.970 ;
        RECT 292.750 245.720 293.290 249.970 ;
        RECT 294.130 245.720 294.670 249.970 ;
        RECT 295.510 245.720 296.050 249.970 ;
        RECT 296.890 245.720 297.430 249.970 ;
        RECT 298.270 245.720 298.810 249.970 ;
        RECT 299.650 245.720 300.190 249.970 ;
        RECT 301.030 245.720 301.570 249.970 ;
        RECT 302.410 245.720 302.950 249.970 ;
        RECT 303.790 245.720 304.330 249.970 ;
        RECT 305.170 245.720 305.710 249.970 ;
        RECT 306.550 245.720 307.090 249.970 ;
        RECT 307.930 245.720 308.470 249.970 ;
        RECT 309.310 245.720 309.850 249.970 ;
        RECT 310.690 245.720 311.230 249.970 ;
        RECT 312.070 245.720 312.610 249.970 ;
        RECT 313.450 245.720 313.990 249.970 ;
        RECT 314.830 245.720 315.370 249.970 ;
        RECT 316.210 245.720 316.750 249.970 ;
        RECT 317.590 245.720 318.130 249.970 ;
        RECT 318.970 245.720 319.510 249.970 ;
        RECT 320.350 245.720 320.890 249.970 ;
        RECT 321.730 245.720 322.270 249.970 ;
        RECT 323.110 245.720 323.650 249.970 ;
        RECT 324.490 245.720 325.030 249.970 ;
        RECT 325.870 245.720 326.410 249.970 ;
        RECT 327.250 245.720 327.790 249.970 ;
        RECT 328.630 245.720 329.170 249.970 ;
        RECT 330.010 245.720 330.550 249.970 ;
        RECT 331.390 245.720 331.930 249.970 ;
        RECT 332.770 245.720 333.310 249.970 ;
        RECT 334.150 245.720 334.690 249.970 ;
        RECT 335.530 245.720 336.070 249.970 ;
        RECT 336.910 245.720 337.450 249.970 ;
        RECT 338.290 245.720 338.830 249.970 ;
        RECT 339.670 245.720 340.210 249.970 ;
        RECT 341.050 245.720 341.590 249.970 ;
        RECT 342.430 245.720 342.970 249.970 ;
        RECT 343.810 245.720 344.350 249.970 ;
        RECT 345.190 245.720 345.730 249.970 ;
        RECT 346.570 245.720 347.110 249.970 ;
        RECT 347.950 245.720 348.490 249.970 ;
        RECT 349.330 245.720 349.870 249.970 ;
        RECT 350.710 245.720 351.250 249.970 ;
        RECT 352.090 245.720 352.630 249.970 ;
        RECT 353.470 245.720 354.010 249.970 ;
        RECT 354.850 245.720 355.390 249.970 ;
        RECT 356.230 245.720 356.770 249.970 ;
        RECT 357.610 245.720 358.150 249.970 ;
        RECT 358.990 245.720 359.530 249.970 ;
        RECT 360.370 245.720 360.910 249.970 ;
        RECT 361.750 245.720 362.290 249.970 ;
        RECT 363.130 245.720 363.670 249.970 ;
        RECT 364.510 245.720 365.050 249.970 ;
        RECT 365.890 245.720 366.430 249.970 ;
        RECT 367.270 245.720 367.810 249.970 ;
        RECT 368.650 245.720 369.190 249.970 ;
        RECT 370.030 245.720 370.570 249.970 ;
        RECT 371.410 245.720 371.950 249.970 ;
        RECT 372.790 245.720 373.330 249.970 ;
        RECT 374.170 245.720 374.710 249.970 ;
        RECT 375.550 245.720 376.090 249.970 ;
        RECT 376.930 245.720 377.470 249.970 ;
        RECT 378.310 245.720 378.850 249.970 ;
        RECT 379.690 245.720 380.230 249.970 ;
        RECT 381.070 245.720 381.610 249.970 ;
        RECT 382.450 245.720 382.990 249.970 ;
        RECT 383.830 245.720 384.370 249.970 ;
        RECT 385.210 245.720 385.750 249.970 ;
        RECT 386.590 245.720 387.130 249.970 ;
        RECT 387.970 245.720 388.510 249.970 ;
        RECT 389.350 245.720 389.890 249.970 ;
        RECT 390.730 245.720 391.270 249.970 ;
        RECT 392.110 245.720 392.650 249.970 ;
        RECT 393.490 245.720 394.030 249.970 ;
        RECT 394.870 245.720 395.410 249.970 ;
        RECT 396.250 245.720 396.790 249.970 ;
        RECT 397.630 245.720 398.170 249.970 ;
        RECT 399.010 245.720 399.550 249.970 ;
        RECT 400.390 245.720 400.930 249.970 ;
        RECT 401.770 245.720 402.310 249.970 ;
        RECT 403.150 245.720 403.690 249.970 ;
        RECT 404.530 245.720 405.070 249.970 ;
        RECT 405.910 245.720 406.450 249.970 ;
        RECT 407.290 245.720 407.830 249.970 ;
        RECT 408.670 245.720 409.210 249.970 ;
        RECT 410.050 245.720 410.590 249.970 ;
        RECT 411.430 245.720 411.970 249.970 ;
        RECT 412.810 245.720 413.350 249.970 ;
        RECT 414.190 245.720 414.730 249.970 ;
        RECT 415.570 245.720 416.110 249.970 ;
        RECT 416.950 245.720 417.490 249.970 ;
        RECT 418.330 245.720 418.870 249.970 ;
        RECT 419.710 245.720 420.250 249.970 ;
        RECT 421.090 245.720 421.630 249.970 ;
        RECT 422.470 245.720 423.010 249.970 ;
        RECT 423.850 245.720 424.390 249.970 ;
        RECT 425.230 245.720 425.770 249.970 ;
        RECT 426.610 245.720 427.150 249.970 ;
        RECT 427.990 245.720 428.530 249.970 ;
        RECT 429.370 245.720 429.910 249.970 ;
        RECT 430.750 245.720 431.290 249.970 ;
        RECT 432.130 245.720 432.670 249.970 ;
        RECT 433.510 245.720 434.050 249.970 ;
        RECT 434.890 245.720 435.430 249.970 ;
        RECT 436.270 245.720 436.810 249.970 ;
        RECT 437.650 245.720 438.190 249.970 ;
        RECT 439.030 245.720 439.570 249.970 ;
        RECT 440.410 245.720 440.950 249.970 ;
        RECT 441.790 245.720 442.330 249.970 ;
        RECT 443.170 245.720 443.710 249.970 ;
        RECT 444.550 245.720 445.090 249.970 ;
        RECT 445.930 245.720 446.470 249.970 ;
        RECT 447.310 245.720 447.850 249.970 ;
        RECT 448.690 245.720 449.230 249.970 ;
        RECT 450.070 245.720 450.610 249.970 ;
        RECT 451.450 245.720 451.990 249.970 ;
        RECT 452.830 245.720 453.370 249.970 ;
        RECT 454.210 245.720 454.750 249.970 ;
        RECT 455.590 245.720 456.130 249.970 ;
        RECT 456.970 245.720 457.510 249.970 ;
        RECT 458.350 245.720 458.890 249.970 ;
        RECT 459.730 245.720 460.270 249.970 ;
        RECT 461.110 245.720 461.650 249.970 ;
        RECT 462.490 245.720 463.030 249.970 ;
        RECT 463.870 245.720 464.410 249.970 ;
        RECT 465.250 245.720 465.790 249.970 ;
        RECT 466.630 245.720 467.170 249.970 ;
        RECT 468.010 245.720 468.550 249.970 ;
        RECT 469.390 245.720 469.930 249.970 ;
        RECT 470.770 245.720 471.310 249.970 ;
        RECT 472.150 245.720 472.690 249.970 ;
        RECT 473.530 245.720 474.070 249.970 ;
        RECT 474.910 245.720 475.450 249.970 ;
        RECT 476.290 245.720 476.830 249.970 ;
        RECT 477.670 245.720 478.210 249.970 ;
        RECT 479.050 245.720 479.590 249.970 ;
        RECT 480.430 245.720 480.970 249.970 ;
        RECT 481.810 245.720 482.350 249.970 ;
        RECT 483.190 245.720 483.730 249.970 ;
        RECT 484.570 245.720 485.110 249.970 ;
        RECT 485.950 245.720 486.490 249.970 ;
        RECT 487.330 245.720 487.870 249.970 ;
        RECT 488.710 245.720 489.250 249.970 ;
        RECT 490.090 245.720 490.630 249.970 ;
        RECT 491.470 245.720 492.010 249.970 ;
        RECT 492.850 245.720 493.390 249.970 ;
        RECT 494.230 245.720 494.770 249.970 ;
        RECT 495.610 245.720 496.150 249.970 ;
        RECT 496.990 245.720 497.530 249.970 ;
        RECT 498.370 245.720 498.910 249.970 ;
        RECT 499.750 245.720 500.290 249.970 ;
        RECT 501.130 245.720 501.670 249.970 ;
        RECT 502.510 245.720 503.050 249.970 ;
        RECT 503.890 245.720 504.430 249.970 ;
        RECT 505.270 245.720 505.810 249.970 ;
        RECT 506.650 245.720 507.190 249.970 ;
        RECT 508.030 245.720 508.570 249.970 ;
        RECT 509.410 245.720 509.950 249.970 ;
        RECT 510.790 245.720 511.330 249.970 ;
        RECT 512.170 245.720 512.710 249.970 ;
        RECT 513.550 245.720 514.090 249.970 ;
        RECT 514.930 245.720 515.470 249.970 ;
        RECT 516.310 245.720 516.850 249.970 ;
        RECT 517.690 245.720 518.230 249.970 ;
        RECT 519.070 245.720 519.610 249.970 ;
        RECT 520.450 245.720 520.990 249.970 ;
        RECT 521.830 245.720 522.370 249.970 ;
        RECT 523.210 245.720 523.750 249.970 ;
        RECT 524.590 245.720 525.130 249.970 ;
        RECT 525.970 245.720 526.510 249.970 ;
        RECT 527.350 245.720 527.890 249.970 ;
        RECT 528.730 245.720 529.270 249.970 ;
        RECT 530.110 245.720 530.650 249.970 ;
        RECT 531.490 245.720 532.030 249.970 ;
        RECT 532.870 245.720 533.410 249.970 ;
        RECT 534.250 245.720 534.790 249.970 ;
        RECT 535.630 245.720 536.170 249.970 ;
        RECT 537.010 245.720 537.550 249.970 ;
        RECT 538.390 245.720 538.930 249.970 ;
        RECT 539.770 245.720 540.310 249.970 ;
        RECT 541.150 245.720 541.690 249.970 ;
        RECT 542.530 245.720 543.070 249.970 ;
        RECT 543.910 245.720 544.450 249.970 ;
        RECT 545.290 245.720 545.830 249.970 ;
        RECT 546.670 245.720 547.210 249.970 ;
        RECT 548.050 245.720 548.590 249.970 ;
        RECT 549.430 245.720 549.970 249.970 ;
        RECT 550.810 245.720 551.350 249.970 ;
        RECT 552.190 245.720 552.730 249.970 ;
        RECT 553.570 245.720 554.110 249.970 ;
        RECT 554.950 245.720 555.490 249.970 ;
        RECT 556.330 245.720 556.870 249.970 ;
        RECT 557.710 245.720 558.250 249.970 ;
        RECT 559.090 245.720 559.630 249.970 ;
        RECT 560.470 245.720 561.010 249.970 ;
        RECT 561.850 245.720 562.390 249.970 ;
        RECT 563.230 245.720 563.770 249.970 ;
        RECT 564.610 245.720 565.150 249.970 ;
        RECT 565.990 245.720 566.530 249.970 ;
        RECT 567.370 245.720 567.910 249.970 ;
        RECT 568.750 245.720 569.290 249.970 ;
        RECT 570.130 245.720 570.670 249.970 ;
        RECT 571.510 245.720 572.050 249.970 ;
        RECT 572.890 245.720 573.430 249.970 ;
        RECT 574.270 245.720 574.810 249.970 ;
        RECT 575.650 245.720 576.190 249.970 ;
        RECT 577.030 245.720 577.570 249.970 ;
        RECT 578.410 245.720 578.950 249.970 ;
        RECT 579.790 245.720 580.330 249.970 ;
        RECT 581.170 245.720 581.710 249.970 ;
        RECT 582.550 245.720 583.090 249.970 ;
        RECT 583.930 245.720 584.470 249.970 ;
        RECT 585.310 245.720 585.850 249.970 ;
        RECT 586.690 245.720 587.230 249.970 ;
        RECT 588.070 245.720 588.610 249.970 ;
        RECT 589.450 245.720 589.990 249.970 ;
        RECT 590.830 245.720 591.370 249.970 ;
        RECT 592.210 245.720 592.750 249.970 ;
        RECT 593.590 245.720 594.130 249.970 ;
        RECT 594.970 245.720 595.510 249.970 ;
        RECT 596.350 245.720 596.890 249.970 ;
        RECT 597.730 245.720 598.270 249.970 ;
        RECT 599.110 245.720 599.650 249.970 ;
        RECT 600.490 245.720 601.030 249.970 ;
        RECT 601.870 245.720 602.410 249.970 ;
        RECT 603.250 245.720 603.790 249.970 ;
        RECT 604.630 245.720 605.170 249.970 ;
        RECT 606.010 245.720 606.550 249.970 ;
        RECT 607.390 245.720 607.930 249.970 ;
        RECT 608.770 245.720 609.310 249.970 ;
        RECT 610.150 245.720 610.690 249.970 ;
        RECT 611.530 245.720 612.070 249.970 ;
        RECT 612.910 245.720 613.450 249.970 ;
        RECT 614.290 245.720 614.830 249.970 ;
        RECT 615.670 245.720 616.210 249.970 ;
        RECT 617.050 245.720 617.590 249.970 ;
        RECT 618.430 245.720 618.970 249.970 ;
        RECT 619.810 245.720 620.350 249.970 ;
        RECT 621.190 245.720 621.730 249.970 ;
        RECT 622.570 245.720 623.110 249.970 ;
        RECT 623.950 245.720 624.490 249.970 ;
        RECT 625.330 245.720 625.870 249.970 ;
        RECT 626.710 245.720 627.250 249.970 ;
        RECT 628.090 245.720 628.630 249.970 ;
        RECT 629.470 245.720 638.380 249.970 ;
        RECT 7.970 4.280 638.380 245.720 ;
        RECT 7.970 4.000 18.670 4.280 ;
        RECT 19.510 4.000 27.410 4.280 ;
        RECT 28.250 4.000 36.150 4.280 ;
        RECT 36.990 4.000 44.890 4.280 ;
        RECT 45.730 4.000 53.630 4.280 ;
        RECT 54.470 4.000 62.370 4.280 ;
        RECT 63.210 4.000 71.110 4.280 ;
        RECT 71.950 4.000 79.850 4.280 ;
        RECT 80.690 4.000 88.590 4.280 ;
        RECT 89.430 4.000 97.330 4.280 ;
        RECT 98.170 4.000 106.070 4.280 ;
        RECT 106.910 4.000 114.810 4.280 ;
        RECT 115.650 4.000 123.550 4.280 ;
        RECT 124.390 4.000 132.290 4.280 ;
        RECT 133.130 4.000 141.030 4.280 ;
        RECT 141.870 4.000 149.770 4.280 ;
        RECT 150.610 4.000 158.510 4.280 ;
        RECT 159.350 4.000 167.250 4.280 ;
        RECT 168.090 4.000 175.990 4.280 ;
        RECT 176.830 4.000 184.730 4.280 ;
        RECT 185.570 4.000 193.470 4.280 ;
        RECT 194.310 4.000 202.210 4.280 ;
        RECT 203.050 4.000 210.950 4.280 ;
        RECT 211.790 4.000 219.690 4.280 ;
        RECT 220.530 4.000 228.430 4.280 ;
        RECT 229.270 4.000 237.170 4.280 ;
        RECT 238.010 4.000 245.910 4.280 ;
        RECT 246.750 4.000 254.650 4.280 ;
        RECT 255.490 4.000 263.390 4.280 ;
        RECT 264.230 4.000 272.130 4.280 ;
        RECT 272.970 4.000 280.870 4.280 ;
        RECT 281.710 4.000 289.610 4.280 ;
        RECT 290.450 4.000 298.350 4.280 ;
        RECT 299.190 4.000 307.090 4.280 ;
        RECT 307.930 4.000 315.830 4.280 ;
        RECT 316.670 4.000 324.570 4.280 ;
        RECT 325.410 4.000 333.310 4.280 ;
        RECT 334.150 4.000 342.050 4.280 ;
        RECT 342.890 4.000 350.790 4.280 ;
        RECT 351.630 4.000 359.530 4.280 ;
        RECT 360.370 4.000 368.270 4.280 ;
        RECT 369.110 4.000 377.010 4.280 ;
        RECT 377.850 4.000 385.750 4.280 ;
        RECT 386.590 4.000 394.490 4.280 ;
        RECT 395.330 4.000 403.230 4.280 ;
        RECT 404.070 4.000 411.970 4.280 ;
        RECT 412.810 4.000 420.710 4.280 ;
        RECT 421.550 4.000 429.450 4.280 ;
        RECT 430.290 4.000 438.190 4.280 ;
        RECT 439.030 4.000 446.930 4.280 ;
        RECT 447.770 4.000 455.670 4.280 ;
        RECT 456.510 4.000 464.410 4.280 ;
        RECT 465.250 4.000 473.150 4.280 ;
        RECT 473.990 4.000 481.890 4.280 ;
        RECT 482.730 4.000 490.630 4.280 ;
        RECT 491.470 4.000 499.370 4.280 ;
        RECT 500.210 4.000 508.110 4.280 ;
        RECT 508.950 4.000 516.850 4.280 ;
        RECT 517.690 4.000 525.590 4.280 ;
        RECT 526.430 4.000 534.330 4.280 ;
        RECT 535.170 4.000 543.070 4.280 ;
        RECT 543.910 4.000 551.810 4.280 ;
        RECT 552.650 4.000 560.550 4.280 ;
        RECT 561.390 4.000 569.290 4.280 ;
        RECT 570.130 4.000 578.030 4.280 ;
        RECT 578.870 4.000 586.770 4.280 ;
        RECT 587.610 4.000 595.510 4.280 ;
        RECT 596.350 4.000 604.250 4.280 ;
        RECT 605.090 4.000 612.990 4.280 ;
        RECT 613.830 4.000 621.730 4.280 ;
        RECT 622.570 4.000 630.470 4.280 ;
        RECT 631.310 4.000 638.380 4.280 ;
      LAYER met3 ;
        RECT 7.950 10.715 637.030 249.385 ;
      LAYER met4 ;
        RECT 19.615 237.280 617.025 245.985 ;
        RECT 19.615 178.760 20.640 237.280 ;
        RECT 23.040 178.760 97.440 237.280 ;
        RECT 99.840 178.760 174.240 237.280 ;
        RECT 176.640 178.760 251.040 237.280 ;
        RECT 253.440 178.760 327.840 237.280 ;
        RECT 330.240 178.760 404.640 237.280 ;
        RECT 407.040 178.760 481.440 237.280 ;
        RECT 483.840 178.760 558.240 237.280 ;
        RECT 560.640 178.760 617.025 237.280 ;
        RECT 19.615 27.480 617.025 178.760 ;
  END
END InstructionCache
END LIBRARY

