VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM32_1RW1R
  CLASS BLOCK ;
  FOREIGN RAM32_1RW1R ;
  ORIGIN 0.000 0.000 ;
  SIZE 592.020 BY 144.160 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 590.020 78.920 592.020 79.520 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 590.020 93.200 592.020 93.800 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 590.020 107.480 592.020 108.080 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 590.020 121.760 592.020 122.360 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 590.020 136.040 592.020 136.640 ;
    END
  END A0[4]
  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 2.000 31.240 ;
    END
  END A1[0]
  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 2.000 51.640 ;
    END
  END A1[1]
  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 2.000 72.040 ;
    END
  END A1[2]
  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 2.000 92.440 ;
    END
  END A1[3]
  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 2.000 112.840 ;
    END
  END A1[4]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 2.000 10.840 ;
    END
  END CLK
  PIN Di0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 0.000 10.950 2.000 ;
    END
  END Di0[0]
  PIN Di0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 0.000 194.950 2.000 ;
    END
  END Di0[10]
  PIN Di0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.070 0.000 213.350 2.000 ;
    END
  END Di0[11]
  PIN Di0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.470 0.000 231.750 2.000 ;
    END
  END Di0[12]
  PIN Di0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 0.000 250.150 2.000 ;
    END
  END Di0[13]
  PIN Di0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 0.000 268.550 2.000 ;
    END
  END Di0[14]
  PIN Di0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 2.000 ;
    END
  END Di0[15]
  PIN Di0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 0.000 305.350 2.000 ;
    END
  END Di0[16]
  PIN Di0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.470 0.000 323.750 2.000 ;
    END
  END Di0[17]
  PIN Di0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.870 0.000 342.150 2.000 ;
    END
  END Di0[18]
  PIN Di0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.270 0.000 360.550 2.000 ;
    END
  END Di0[19]
  PIN Di0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 2.000 ;
    END
  END Di0[1]
  PIN Di0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.670 0.000 378.950 2.000 ;
    END
  END Di0[20]
  PIN Di0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.070 0.000 397.350 2.000 ;
    END
  END Di0[21]
  PIN Di0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 0.000 415.750 2.000 ;
    END
  END Di0[22]
  PIN Di0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.870 0.000 434.150 2.000 ;
    END
  END Di0[23]
  PIN Di0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.270 0.000 452.550 2.000 ;
    END
  END Di0[24]
  PIN Di0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.670 0.000 470.950 2.000 ;
    END
  END Di0[25]
  PIN Di0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.070 0.000 489.350 2.000 ;
    END
  END Di0[26]
  PIN Di0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.470 0.000 507.750 2.000 ;
    END
  END Di0[27]
  PIN Di0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.870 0.000 526.150 2.000 ;
    END
  END Di0[28]
  PIN Di0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 0.000 544.550 2.000 ;
    END
  END Di0[29]
  PIN Di0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 0.000 47.750 2.000 ;
    END
  END Di0[2]
  PIN Di0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.670 0.000 562.950 2.000 ;
    END
  END Di0[30]
  PIN Di0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.070 0.000 581.350 2.000 ;
    END
  END Di0[31]
  PIN Di0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 0.000 66.150 2.000 ;
    END
  END Di0[3]
  PIN Di0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 0.000 84.550 2.000 ;
    END
  END Di0[4]
  PIN Di0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 0.000 102.950 2.000 ;
    END
  END Di0[5]
  PIN Di0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.070 0.000 121.350 2.000 ;
    END
  END Di0[6]
  PIN Di0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 0.000 139.750 2.000 ;
    END
  END Di0[7]
  PIN Di0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 2.000 ;
    END
  END Di0[8]
  PIN Di0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 0.000 176.550 2.000 ;
    END
  END Di0[9]
  PIN Do0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 142.160 6.350 144.160 ;
    END
  END Do0[0]
  PIN Do0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 142.160 98.350 144.160 ;
    END
  END Do0[10]
  PIN Do0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 142.160 116.750 144.160 ;
    END
  END Do0[11]
  PIN Do0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.870 142.160 135.150 144.160 ;
    END
  END Do0[12]
  PIN Do0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 142.160 153.550 144.160 ;
    END
  END Do0[13]
  PIN Do0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 142.160 171.950 144.160 ;
    END
  END Do0[14]
  PIN Do0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 142.160 190.350 144.160 ;
    END
  END Do0[15]
  PIN Do0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 142.160 208.750 144.160 ;
    END
  END Do0[16]
  PIN Do0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.870 142.160 227.150 144.160 ;
    END
  END Do0[17]
  PIN Do0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.270 142.160 245.550 144.160 ;
    END
  END Do0[18]
  PIN Do0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 142.160 263.950 144.160 ;
    END
  END Do0[19]
  PIN Do0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 142.160 15.550 144.160 ;
    END
  END Do0[1]
  PIN Do0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.070 142.160 282.350 144.160 ;
    END
  END Do0[20]
  PIN Do0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.270 142.160 291.550 144.160 ;
    END
  END Do0[21]
  PIN Do0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.470 142.160 300.750 144.160 ;
    END
  END Do0[22]
  PIN Do0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.670 142.160 309.950 144.160 ;
    END
  END Do0[23]
  PIN Do0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 142.160 319.150 144.160 ;
    END
  END Do0[24]
  PIN Do0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.070 142.160 328.350 144.160 ;
    END
  END Do0[25]
  PIN Do0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.270 142.160 337.550 144.160 ;
    END
  END Do0[26]
  PIN Do0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.470 142.160 346.750 144.160 ;
    END
  END Do0[27]
  PIN Do0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.670 142.160 355.950 144.160 ;
    END
  END Do0[28]
  PIN Do0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.870 142.160 365.150 144.160 ;
    END
  END Do0[29]
  PIN Do0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 142.160 24.750 144.160 ;
    END
  END Do0[2]
  PIN Do0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.070 142.160 374.350 144.160 ;
    END
  END Do0[30]
  PIN Do0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 142.160 383.550 144.160 ;
    END
  END Do0[31]
  PIN Do0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 142.160 33.950 144.160 ;
    END
  END Do0[3]
  PIN Do0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 142.160 43.150 144.160 ;
    END
  END Do0[4]
  PIN Do0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 142.160 52.350 144.160 ;
    END
  END Do0[5]
  PIN Do0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 142.160 61.550 144.160 ;
    END
  END Do0[6]
  PIN Do0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 142.160 70.750 144.160 ;
    END
  END Do0[7]
  PIN Do0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 142.160 79.950 144.160 ;
    END
  END Do0[8]
  PIN Do0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 142.160 89.150 144.160 ;
    END
  END Do0[9]
  PIN Do1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 142.160 107.550 144.160 ;
    END
  END Do1[0]
  PIN Do1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.470 142.160 392.750 144.160 ;
    END
  END Do1[10]
  PIN Do1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.670 142.160 401.950 144.160 ;
    END
  END Do1[11]
  PIN Do1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.870 142.160 411.150 144.160 ;
    END
  END Do1[12]
  PIN Do1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.070 142.160 420.350 144.160 ;
    END
  END Do1[13]
  PIN Do1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.270 142.160 429.550 144.160 ;
    END
  END Do1[14]
  PIN Do1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.470 142.160 438.750 144.160 ;
    END
  END Do1[15]
  PIN Do1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 142.160 447.950 144.160 ;
    END
  END Do1[16]
  PIN Do1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.870 142.160 457.150 144.160 ;
    END
  END Do1[17]
  PIN Do1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.070 142.160 466.350 144.160 ;
    END
  END Do1[18]
  PIN Do1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.270 142.160 475.550 144.160 ;
    END
  END Do1[19]
  PIN Do1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 142.160 125.950 144.160 ;
    END
  END Do1[1]
  PIN Do1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.470 142.160 484.750 144.160 ;
    END
  END Do1[20]
  PIN Do1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.670 142.160 493.950 144.160 ;
    END
  END Do1[21]
  PIN Do1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.870 142.160 503.150 144.160 ;
    END
  END Do1[22]
  PIN Do1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 142.160 512.350 144.160 ;
    END
  END Do1[23]
  PIN Do1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.270 142.160 521.550 144.160 ;
    END
  END Do1[24]
  PIN Do1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.470 142.160 530.750 144.160 ;
    END
  END Do1[25]
  PIN Do1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.670 142.160 539.950 144.160 ;
    END
  END Do1[26]
  PIN Do1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.870 142.160 549.150 144.160 ;
    END
  END Do1[27]
  PIN Do1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.070 142.160 558.350 144.160 ;
    END
  END Do1[28]
  PIN Do1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.270 142.160 567.550 144.160 ;
    END
  END Do1[29]
  PIN Do1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 142.160 144.350 144.160 ;
    END
  END Do1[2]
  PIN Do1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.470 142.160 576.750 144.160 ;
    END
  END Do1[30]
  PIN Do1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.670 142.160 585.950 144.160 ;
    END
  END Do1[31]
  PIN Do1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.470 142.160 162.750 144.160 ;
    END
  END Do1[3]
  PIN Do1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.870 142.160 181.150 144.160 ;
    END
  END Do1[4]
  PIN Do1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.270 142.160 199.550 144.160 ;
    END
  END Do1[5]
  PIN Do1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 142.160 217.950 144.160 ;
    END
  END Do1[6]
  PIN Do1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 142.160 236.350 144.160 ;
    END
  END Do1[7]
  PIN Do1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 142.160 254.750 144.160 ;
    END
  END Do1[8]
  PIN Do1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.870 142.160 273.150 144.160 ;
    END
  END Do1[9]
  PIN EN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 590.020 7.520 592.020 8.120 ;
    END
  END EN0
  PIN EN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 2.000 133.240 ;
    END
  END EN1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 95.080 2.480 96.680 141.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 248.680 2.480 250.280 141.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 402.280 2.480 403.880 141.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 555.880 2.480 557.480 141.680 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 18.280 2.480 19.880 141.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.880 2.480 173.480 141.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.480 2.480 327.080 141.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 479.080 2.480 480.680 141.680 ;
    END
  END VPWR
  PIN WE0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 590.020 21.800 592.020 22.400 ;
    END
  END WE0[0]
  PIN WE0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 590.020 36.080 592.020 36.680 ;
    END
  END WE0[1]
  PIN WE0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 590.020 50.360 592.020 50.960 ;
    END
  END WE0[2]
  PIN WE0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 590.020 64.640 592.020 65.240 ;
    END
  END WE0[3]
  OBS
      LAYER li1 ;
        RECT 2.760 2.635 589.260 141.525 ;
      LAYER met1 ;
        RECT 1.450 0.040 589.260 144.120 ;
      LAYER met2 ;
        RECT 1.480 141.880 5.790 144.150 ;
        RECT 6.630 141.880 14.990 144.150 ;
        RECT 15.830 141.880 24.190 144.150 ;
        RECT 25.030 141.880 33.390 144.150 ;
        RECT 34.230 141.880 42.590 144.150 ;
        RECT 43.430 141.880 51.790 144.150 ;
        RECT 52.630 141.880 60.990 144.150 ;
        RECT 61.830 141.880 70.190 144.150 ;
        RECT 71.030 141.880 79.390 144.150 ;
        RECT 80.230 141.880 88.590 144.150 ;
        RECT 89.430 141.880 97.790 144.150 ;
        RECT 98.630 141.880 106.990 144.150 ;
        RECT 107.830 141.880 116.190 144.150 ;
        RECT 117.030 141.880 125.390 144.150 ;
        RECT 126.230 141.880 134.590 144.150 ;
        RECT 135.430 141.880 143.790 144.150 ;
        RECT 144.630 141.880 152.990 144.150 ;
        RECT 153.830 141.880 162.190 144.150 ;
        RECT 163.030 141.880 171.390 144.150 ;
        RECT 172.230 141.880 180.590 144.150 ;
        RECT 181.430 141.880 189.790 144.150 ;
        RECT 190.630 141.880 198.990 144.150 ;
        RECT 199.830 141.880 208.190 144.150 ;
        RECT 209.030 141.880 217.390 144.150 ;
        RECT 218.230 141.880 226.590 144.150 ;
        RECT 227.430 141.880 235.790 144.150 ;
        RECT 236.630 141.880 244.990 144.150 ;
        RECT 245.830 141.880 254.190 144.150 ;
        RECT 255.030 141.880 263.390 144.150 ;
        RECT 264.230 141.880 272.590 144.150 ;
        RECT 273.430 141.880 281.790 144.150 ;
        RECT 282.630 141.880 290.990 144.150 ;
        RECT 291.830 141.880 300.190 144.150 ;
        RECT 301.030 141.880 309.390 144.150 ;
        RECT 310.230 141.880 318.590 144.150 ;
        RECT 319.430 141.880 327.790 144.150 ;
        RECT 328.630 141.880 336.990 144.150 ;
        RECT 337.830 141.880 346.190 144.150 ;
        RECT 347.030 141.880 355.390 144.150 ;
        RECT 356.230 141.880 364.590 144.150 ;
        RECT 365.430 141.880 373.790 144.150 ;
        RECT 374.630 141.880 382.990 144.150 ;
        RECT 383.830 141.880 392.190 144.150 ;
        RECT 393.030 141.880 401.390 144.150 ;
        RECT 402.230 141.880 410.590 144.150 ;
        RECT 411.430 141.880 419.790 144.150 ;
        RECT 420.630 141.880 428.990 144.150 ;
        RECT 429.830 141.880 438.190 144.150 ;
        RECT 439.030 141.880 447.390 144.150 ;
        RECT 448.230 141.880 456.590 144.150 ;
        RECT 457.430 141.880 465.790 144.150 ;
        RECT 466.630 141.880 474.990 144.150 ;
        RECT 475.830 141.880 484.190 144.150 ;
        RECT 485.030 141.880 493.390 144.150 ;
        RECT 494.230 141.880 502.590 144.150 ;
        RECT 503.430 141.880 511.790 144.150 ;
        RECT 512.630 141.880 520.990 144.150 ;
        RECT 521.830 141.880 530.190 144.150 ;
        RECT 531.030 141.880 539.390 144.150 ;
        RECT 540.230 141.880 548.590 144.150 ;
        RECT 549.430 141.880 557.790 144.150 ;
        RECT 558.630 141.880 566.990 144.150 ;
        RECT 567.830 141.880 576.190 144.150 ;
        RECT 577.030 141.880 585.390 144.150 ;
        RECT 1.480 2.280 585.940 141.880 ;
        RECT 1.480 0.010 10.390 2.280 ;
        RECT 11.230 0.010 28.790 2.280 ;
        RECT 29.630 0.010 47.190 2.280 ;
        RECT 48.030 0.010 65.590 2.280 ;
        RECT 66.430 0.010 83.990 2.280 ;
        RECT 84.830 0.010 102.390 2.280 ;
        RECT 103.230 0.010 120.790 2.280 ;
        RECT 121.630 0.010 139.190 2.280 ;
        RECT 140.030 0.010 157.590 2.280 ;
        RECT 158.430 0.010 175.990 2.280 ;
        RECT 176.830 0.010 194.390 2.280 ;
        RECT 195.230 0.010 212.790 2.280 ;
        RECT 213.630 0.010 231.190 2.280 ;
        RECT 232.030 0.010 249.590 2.280 ;
        RECT 250.430 0.010 267.990 2.280 ;
        RECT 268.830 0.010 286.390 2.280 ;
        RECT 287.230 0.010 304.790 2.280 ;
        RECT 305.630 0.010 323.190 2.280 ;
        RECT 324.030 0.010 341.590 2.280 ;
        RECT 342.430 0.010 359.990 2.280 ;
        RECT 360.830 0.010 378.390 2.280 ;
        RECT 379.230 0.010 396.790 2.280 ;
        RECT 397.630 0.010 415.190 2.280 ;
        RECT 416.030 0.010 433.590 2.280 ;
        RECT 434.430 0.010 451.990 2.280 ;
        RECT 452.830 0.010 470.390 2.280 ;
        RECT 471.230 0.010 488.790 2.280 ;
        RECT 489.630 0.010 507.190 2.280 ;
        RECT 508.030 0.010 525.590 2.280 ;
        RECT 526.430 0.010 543.990 2.280 ;
        RECT 544.830 0.010 562.390 2.280 ;
        RECT 563.230 0.010 580.790 2.280 ;
        RECT 581.630 0.010 585.940 2.280 ;
      LAYER met3 ;
        RECT 2.000 137.040 590.020 143.305 ;
        RECT 2.000 135.640 589.620 137.040 ;
        RECT 2.000 133.640 590.020 135.640 ;
        RECT 2.400 132.240 590.020 133.640 ;
        RECT 2.000 122.760 590.020 132.240 ;
        RECT 2.000 121.360 589.620 122.760 ;
        RECT 2.000 113.240 590.020 121.360 ;
        RECT 2.400 111.840 590.020 113.240 ;
        RECT 2.000 108.480 590.020 111.840 ;
        RECT 2.000 107.080 589.620 108.480 ;
        RECT 2.000 94.200 590.020 107.080 ;
        RECT 2.000 92.840 589.620 94.200 ;
        RECT 2.400 92.800 589.620 92.840 ;
        RECT 2.400 91.440 590.020 92.800 ;
        RECT 2.000 79.920 590.020 91.440 ;
        RECT 2.000 78.520 589.620 79.920 ;
        RECT 2.000 72.440 590.020 78.520 ;
        RECT 2.400 71.040 590.020 72.440 ;
        RECT 2.000 65.640 590.020 71.040 ;
        RECT 2.000 64.240 589.620 65.640 ;
        RECT 2.000 52.040 590.020 64.240 ;
        RECT 2.400 51.360 590.020 52.040 ;
        RECT 2.400 50.640 589.620 51.360 ;
        RECT 2.000 49.960 589.620 50.640 ;
        RECT 2.000 37.080 590.020 49.960 ;
        RECT 2.000 35.680 589.620 37.080 ;
        RECT 2.000 31.640 590.020 35.680 ;
        RECT 2.400 30.240 590.020 31.640 ;
        RECT 2.000 22.800 590.020 30.240 ;
        RECT 2.000 21.400 589.620 22.800 ;
        RECT 2.000 11.240 590.020 21.400 ;
        RECT 2.400 9.840 590.020 11.240 ;
        RECT 2.000 8.520 590.020 9.840 ;
        RECT 2.000 7.120 589.620 8.520 ;
        RECT 2.000 0.175 590.020 7.120 ;
      LAYER met4 ;
        RECT 8.575 13.095 17.880 126.985 ;
        RECT 20.280 13.095 94.680 126.985 ;
        RECT 97.080 13.095 171.480 126.985 ;
        RECT 173.880 13.095 248.280 126.985 ;
        RECT 250.680 13.095 325.080 126.985 ;
        RECT 327.480 13.095 401.880 126.985 ;
        RECT 404.280 13.095 478.680 126.985 ;
        RECT 481.080 13.095 544.345 126.985 ;
  END
END RAM32_1RW1R
END LIBRARY

