module SEL_32x3 (
  input      [31:0]   src0,
  input      [31:0]   src1,
  input      [31:0]   src2,
  input      [2:0]    sel,
  output reg [31:0]   result
);
endmodule