VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DataCache
  CLASS BLOCK ;
  FOREIGN DataCache ;
  ORIGIN 0.000 0.000 ;
  SIZE 650.000 BY 250.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 600.850 246.000 601.130 250.000 ;
    END
  END clk
  PIN io_cpu_execute_address[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 246.000 100.650 250.000 ;
    END
  END io_cpu_execute_address[0]
  PIN io_cpu_execute_address[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 246.000 277.290 250.000 ;
    END
  END io_cpu_execute_address[10]
  PIN io_cpu_execute_address[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.730 246.000 292.010 250.000 ;
    END
  END io_cpu_execute_address[11]
  PIN io_cpu_execute_address[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 246.000 306.730 250.000 ;
    END
  END io_cpu_execute_address[12]
  PIN io_cpu_execute_address[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.170 246.000 321.450 250.000 ;
    END
  END io_cpu_execute_address[13]
  PIN io_cpu_execute_address[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.890 246.000 336.170 250.000 ;
    END
  END io_cpu_execute_address[14]
  PIN io_cpu_execute_address[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.610 246.000 350.890 250.000 ;
    END
  END io_cpu_execute_address[15]
  PIN io_cpu_execute_address[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.330 246.000 365.610 250.000 ;
    END
  END io_cpu_execute_address[16]
  PIN io_cpu_execute_address[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 246.000 380.330 250.000 ;
    END
  END io_cpu_execute_address[17]
  PIN io_cpu_execute_address[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.770 246.000 395.050 250.000 ;
    END
  END io_cpu_execute_address[18]
  PIN io_cpu_execute_address[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.490 246.000 409.770 250.000 ;
    END
  END io_cpu_execute_address[19]
  PIN io_cpu_execute_address[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 246.000 120.890 250.000 ;
    END
  END io_cpu_execute_address[1]
  PIN io_cpu_execute_address[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.210 246.000 424.490 250.000 ;
    END
  END io_cpu_execute_address[20]
  PIN io_cpu_execute_address[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.930 246.000 439.210 250.000 ;
    END
  END io_cpu_execute_address[21]
  PIN io_cpu_execute_address[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.650 246.000 453.930 250.000 ;
    END
  END io_cpu_execute_address[22]
  PIN io_cpu_execute_address[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.370 246.000 468.650 250.000 ;
    END
  END io_cpu_execute_address[23]
  PIN io_cpu_execute_address[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 246.000 483.370 250.000 ;
    END
  END io_cpu_execute_address[24]
  PIN io_cpu_execute_address[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.810 246.000 498.090 250.000 ;
    END
  END io_cpu_execute_address[25]
  PIN io_cpu_execute_address[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.530 246.000 512.810 250.000 ;
    END
  END io_cpu_execute_address[26]
  PIN io_cpu_execute_address[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.250 246.000 527.530 250.000 ;
    END
  END io_cpu_execute_address[27]
  PIN io_cpu_execute_address[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.970 246.000 542.250 250.000 ;
    END
  END io_cpu_execute_address[28]
  PIN io_cpu_execute_address[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 246.000 556.970 250.000 ;
    END
  END io_cpu_execute_address[29]
  PIN io_cpu_execute_address[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 246.000 141.130 250.000 ;
    END
  END io_cpu_execute_address[2]
  PIN io_cpu_execute_address[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.410 246.000 571.690 250.000 ;
    END
  END io_cpu_execute_address[30]
  PIN io_cpu_execute_address[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.130 246.000 586.410 250.000 ;
    END
  END io_cpu_execute_address[31]
  PIN io_cpu_execute_address[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 246.000 159.530 250.000 ;
    END
  END io_cpu_execute_address[3]
  PIN io_cpu_execute_address[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 246.000 177.930 250.000 ;
    END
  END io_cpu_execute_address[4]
  PIN io_cpu_execute_address[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 246.000 194.490 250.000 ;
    END
  END io_cpu_execute_address[5]
  PIN io_cpu_execute_address[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.770 246.000 211.050 250.000 ;
    END
  END io_cpu_execute_address[6]
  PIN io_cpu_execute_address[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.330 246.000 227.610 250.000 ;
    END
  END io_cpu_execute_address[7]
  PIN io_cpu_execute_address[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.890 246.000 244.170 250.000 ;
    END
  END io_cpu_execute_address[8]
  PIN io_cpu_execute_address[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.450 246.000 260.730 250.000 ;
    END
  END io_cpu_execute_address[9]
  PIN io_cpu_execute_args_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 246.000 102.490 250.000 ;
    END
  END io_cpu_execute_args_data[0]
  PIN io_cpu_execute_args_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.850 246.000 279.130 250.000 ;
    END
  END io_cpu_execute_args_data[10]
  PIN io_cpu_execute_args_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 246.000 293.850 250.000 ;
    END
  END io_cpu_execute_args_data[11]
  PIN io_cpu_execute_args_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 246.000 308.570 250.000 ;
    END
  END io_cpu_execute_args_data[12]
  PIN io_cpu_execute_args_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 246.000 323.290 250.000 ;
    END
  END io_cpu_execute_args_data[13]
  PIN io_cpu_execute_args_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.730 246.000 338.010 250.000 ;
    END
  END io_cpu_execute_args_data[14]
  PIN io_cpu_execute_args_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.450 246.000 352.730 250.000 ;
    END
  END io_cpu_execute_args_data[15]
  PIN io_cpu_execute_args_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 246.000 367.450 250.000 ;
    END
  END io_cpu_execute_args_data[16]
  PIN io_cpu_execute_args_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.890 246.000 382.170 250.000 ;
    END
  END io_cpu_execute_args_data[17]
  PIN io_cpu_execute_args_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.610 246.000 396.890 250.000 ;
    END
  END io_cpu_execute_args_data[18]
  PIN io_cpu_execute_args_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.330 246.000 411.610 250.000 ;
    END
  END io_cpu_execute_args_data[19]
  PIN io_cpu_execute_args_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 246.000 122.730 250.000 ;
    END
  END io_cpu_execute_args_data[1]
  PIN io_cpu_execute_args_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.050 246.000 426.330 250.000 ;
    END
  END io_cpu_execute_args_data[20]
  PIN io_cpu_execute_args_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.770 246.000 441.050 250.000 ;
    END
  END io_cpu_execute_args_data[21]
  PIN io_cpu_execute_args_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.490 246.000 455.770 250.000 ;
    END
  END io_cpu_execute_args_data[22]
  PIN io_cpu_execute_args_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 246.000 470.490 250.000 ;
    END
  END io_cpu_execute_args_data[23]
  PIN io_cpu_execute_args_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.930 246.000 485.210 250.000 ;
    END
  END io_cpu_execute_args_data[24]
  PIN io_cpu_execute_args_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.650 246.000 499.930 250.000 ;
    END
  END io_cpu_execute_args_data[25]
  PIN io_cpu_execute_args_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.370 246.000 514.650 250.000 ;
    END
  END io_cpu_execute_args_data[26]
  PIN io_cpu_execute_args_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.090 246.000 529.370 250.000 ;
    END
  END io_cpu_execute_args_data[27]
  PIN io_cpu_execute_args_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.810 246.000 544.090 250.000 ;
    END
  END io_cpu_execute_args_data[28]
  PIN io_cpu_execute_args_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.530 246.000 558.810 250.000 ;
    END
  END io_cpu_execute_args_data[29]
  PIN io_cpu_execute_args_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 246.000 142.970 250.000 ;
    END
  END io_cpu_execute_args_data[2]
  PIN io_cpu_execute_args_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 246.000 573.530 250.000 ;
    END
  END io_cpu_execute_args_data[30]
  PIN io_cpu_execute_args_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.970 246.000 588.250 250.000 ;
    END
  END io_cpu_execute_args_data[31]
  PIN io_cpu_execute_args_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 246.000 161.370 250.000 ;
    END
  END io_cpu_execute_args_data[3]
  PIN io_cpu_execute_args_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 246.000 179.770 250.000 ;
    END
  END io_cpu_execute_args_data[4]
  PIN io_cpu_execute_args_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.050 246.000 196.330 250.000 ;
    END
  END io_cpu_execute_args_data[5]
  PIN io_cpu_execute_args_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 246.000 212.890 250.000 ;
    END
  END io_cpu_execute_args_data[6]
  PIN io_cpu_execute_args_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.170 246.000 229.450 250.000 ;
    END
  END io_cpu_execute_args_data[7]
  PIN io_cpu_execute_args_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.730 246.000 246.010 250.000 ;
    END
  END io_cpu_execute_args_data[8]
  PIN io_cpu_execute_args_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 246.000 262.570 250.000 ;
    END
  END io_cpu_execute_args_data[9]
  PIN io_cpu_execute_args_size[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 246.000 104.330 250.000 ;
    END
  END io_cpu_execute_args_size[0]
  PIN io_cpu_execute_args_size[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 246.000 124.570 250.000 ;
    END
  END io_cpu_execute_args_size[1]
  PIN io_cpu_execute_args_wr
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 246.000 47.290 250.000 ;
    END
  END io_cpu_execute_args_wr
  PIN io_cpu_execute_isValid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 246.000 49.130 250.000 ;
    END
  END io_cpu_execute_isValid
  PIN io_cpu_flush_ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 246.000 50.970 250.000 ;
    END
  END io_cpu_flush_ready
  PIN io_cpu_flush_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 246.000 52.810 250.000 ;
    END
  END io_cpu_flush_valid
  PIN io_cpu_memory_address[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 246.000 106.170 250.000 ;
    END
  END io_cpu_memory_address[0]
  PIN io_cpu_memory_address[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 246.000 280.970 250.000 ;
    END
  END io_cpu_memory_address[10]
  PIN io_cpu_memory_address[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.410 246.000 295.690 250.000 ;
    END
  END io_cpu_memory_address[11]
  PIN io_cpu_memory_address[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.130 246.000 310.410 250.000 ;
    END
  END io_cpu_memory_address[12]
  PIN io_cpu_memory_address[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.850 246.000 325.130 250.000 ;
    END
  END io_cpu_memory_address[13]
  PIN io_cpu_memory_address[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.570 246.000 339.850 250.000 ;
    END
  END io_cpu_memory_address[14]
  PIN io_cpu_memory_address[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 246.000 354.570 250.000 ;
    END
  END io_cpu_memory_address[15]
  PIN io_cpu_memory_address[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.010 246.000 369.290 250.000 ;
    END
  END io_cpu_memory_address[16]
  PIN io_cpu_memory_address[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.730 246.000 384.010 250.000 ;
    END
  END io_cpu_memory_address[17]
  PIN io_cpu_memory_address[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.450 246.000 398.730 250.000 ;
    END
  END io_cpu_memory_address[18]
  PIN io_cpu_memory_address[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.170 246.000 413.450 250.000 ;
    END
  END io_cpu_memory_address[19]
  PIN io_cpu_memory_address[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 246.000 126.410 250.000 ;
    END
  END io_cpu_memory_address[1]
  PIN io_cpu_memory_address[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.890 246.000 428.170 250.000 ;
    END
  END io_cpu_memory_address[20]
  PIN io_cpu_memory_address[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.610 246.000 442.890 250.000 ;
    END
  END io_cpu_memory_address[21]
  PIN io_cpu_memory_address[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 246.000 457.610 250.000 ;
    END
  END io_cpu_memory_address[22]
  PIN io_cpu_memory_address[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.050 246.000 472.330 250.000 ;
    END
  END io_cpu_memory_address[23]
  PIN io_cpu_memory_address[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.770 246.000 487.050 250.000 ;
    END
  END io_cpu_memory_address[24]
  PIN io_cpu_memory_address[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.490 246.000 501.770 250.000 ;
    END
  END io_cpu_memory_address[25]
  PIN io_cpu_memory_address[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.210 246.000 516.490 250.000 ;
    END
  END io_cpu_memory_address[26]
  PIN io_cpu_memory_address[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.930 246.000 531.210 250.000 ;
    END
  END io_cpu_memory_address[27]
  PIN io_cpu_memory_address[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.650 246.000 545.930 250.000 ;
    END
  END io_cpu_memory_address[28]
  PIN io_cpu_memory_address[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 246.000 560.650 250.000 ;
    END
  END io_cpu_memory_address[29]
  PIN io_cpu_memory_address[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 246.000 144.810 250.000 ;
    END
  END io_cpu_memory_address[2]
  PIN io_cpu_memory_address[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.090 246.000 575.370 250.000 ;
    END
  END io_cpu_memory_address[30]
  PIN io_cpu_memory_address[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.810 246.000 590.090 250.000 ;
    END
  END io_cpu_memory_address[31]
  PIN io_cpu_memory_address[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.930 246.000 163.210 250.000 ;
    END
  END io_cpu_memory_address[3]
  PIN io_cpu_memory_address[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.330 246.000 181.610 250.000 ;
    END
  END io_cpu_memory_address[4]
  PIN io_cpu_memory_address[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 246.000 198.170 250.000 ;
    END
  END io_cpu_memory_address[5]
  PIN io_cpu_memory_address[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 246.000 214.730 250.000 ;
    END
  END io_cpu_memory_address[6]
  PIN io_cpu_memory_address[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 246.000 231.290 250.000 ;
    END
  END io_cpu_memory_address[7]
  PIN io_cpu_memory_address[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.570 246.000 247.850 250.000 ;
    END
  END io_cpu_memory_address[8]
  PIN io_cpu_memory_address[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 246.000 264.410 250.000 ;
    END
  END io_cpu_memory_address[9]
  PIN io_cpu_memory_bypassTranslation
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 246.000 54.650 250.000 ;
    END
  END io_cpu_memory_bypassTranslation
  PIN io_cpu_memory_isRemoved
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 246.000 56.490 250.000 ;
    END
  END io_cpu_memory_isRemoved
  PIN io_cpu_memory_isStuck
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 246.000 58.330 250.000 ;
    END
  END io_cpu_memory_isStuck
  PIN io_cpu_memory_isValid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 246.000 60.170 250.000 ;
    END
  END io_cpu_memory_isValid
  PIN io_cpu_memory_isWrite
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 246.000 62.010 250.000 ;
    END
  END io_cpu_memory_isWrite
  PIN io_cpu_memory_mmuBus_busy
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 246.000 63.850 250.000 ;
    END
  END io_cpu_memory_mmuBus_busy
  PIN io_cpu_memory_mmuBus_cmd_bypassTranslation
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 246.000 65.690 250.000 ;
    END
  END io_cpu_memory_mmuBus_cmd_bypassTranslation
  PIN io_cpu_memory_mmuBus_cmd_isValid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 246.000 67.530 250.000 ;
    END
  END io_cpu_memory_mmuBus_cmd_isValid
  PIN io_cpu_memory_mmuBus_cmd_virtualAddress[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 246.000 108.010 250.000 ;
    END
  END io_cpu_memory_mmuBus_cmd_virtualAddress[0]
  PIN io_cpu_memory_mmuBus_cmd_virtualAddress[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.530 246.000 282.810 250.000 ;
    END
  END io_cpu_memory_mmuBus_cmd_virtualAddress[10]
  PIN io_cpu_memory_mmuBus_cmd_virtualAddress[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 246.000 297.530 250.000 ;
    END
  END io_cpu_memory_mmuBus_cmd_virtualAddress[11]
  PIN io_cpu_memory_mmuBus_cmd_virtualAddress[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 246.000 312.250 250.000 ;
    END
  END io_cpu_memory_mmuBus_cmd_virtualAddress[12]
  PIN io_cpu_memory_mmuBus_cmd_virtualAddress[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 246.000 326.970 250.000 ;
    END
  END io_cpu_memory_mmuBus_cmd_virtualAddress[13]
  PIN io_cpu_memory_mmuBus_cmd_virtualAddress[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 246.000 341.690 250.000 ;
    END
  END io_cpu_memory_mmuBus_cmd_virtualAddress[14]
  PIN io_cpu_memory_mmuBus_cmd_virtualAddress[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.130 246.000 356.410 250.000 ;
    END
  END io_cpu_memory_mmuBus_cmd_virtualAddress[15]
  PIN io_cpu_memory_mmuBus_cmd_virtualAddress[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.850 246.000 371.130 250.000 ;
    END
  END io_cpu_memory_mmuBus_cmd_virtualAddress[16]
  PIN io_cpu_memory_mmuBus_cmd_virtualAddress[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.570 246.000 385.850 250.000 ;
    END
  END io_cpu_memory_mmuBus_cmd_virtualAddress[17]
  PIN io_cpu_memory_mmuBus_cmd_virtualAddress[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.290 246.000 400.570 250.000 ;
    END
  END io_cpu_memory_mmuBus_cmd_virtualAddress[18]
  PIN io_cpu_memory_mmuBus_cmd_virtualAddress[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.010 246.000 415.290 250.000 ;
    END
  END io_cpu_memory_mmuBus_cmd_virtualAddress[19]
  PIN io_cpu_memory_mmuBus_cmd_virtualAddress[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.970 246.000 128.250 250.000 ;
    END
  END io_cpu_memory_mmuBus_cmd_virtualAddress[1]
  PIN io_cpu_memory_mmuBus_cmd_virtualAddress[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.730 246.000 430.010 250.000 ;
    END
  END io_cpu_memory_mmuBus_cmd_virtualAddress[20]
  PIN io_cpu_memory_mmuBus_cmd_virtualAddress[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 246.000 444.730 250.000 ;
    END
  END io_cpu_memory_mmuBus_cmd_virtualAddress[21]
  PIN io_cpu_memory_mmuBus_cmd_virtualAddress[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.170 246.000 459.450 250.000 ;
    END
  END io_cpu_memory_mmuBus_cmd_virtualAddress[22]
  PIN io_cpu_memory_mmuBus_cmd_virtualAddress[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.890 246.000 474.170 250.000 ;
    END
  END io_cpu_memory_mmuBus_cmd_virtualAddress[23]
  PIN io_cpu_memory_mmuBus_cmd_virtualAddress[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.610 246.000 488.890 250.000 ;
    END
  END io_cpu_memory_mmuBus_cmd_virtualAddress[24]
  PIN io_cpu_memory_mmuBus_cmd_virtualAddress[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.330 246.000 503.610 250.000 ;
    END
  END io_cpu_memory_mmuBus_cmd_virtualAddress[25]
  PIN io_cpu_memory_mmuBus_cmd_virtualAddress[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.050 246.000 518.330 250.000 ;
    END
  END io_cpu_memory_mmuBus_cmd_virtualAddress[26]
  PIN io_cpu_memory_mmuBus_cmd_virtualAddress[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.770 246.000 533.050 250.000 ;
    END
  END io_cpu_memory_mmuBus_cmd_virtualAddress[27]
  PIN io_cpu_memory_mmuBus_cmd_virtualAddress[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 246.000 547.770 250.000 ;
    END
  END io_cpu_memory_mmuBus_cmd_virtualAddress[28]
  PIN io_cpu_memory_mmuBus_cmd_virtualAddress[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.210 246.000 562.490 250.000 ;
    END
  END io_cpu_memory_mmuBus_cmd_virtualAddress[29]
  PIN io_cpu_memory_mmuBus_cmd_virtualAddress[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 246.000 146.650 250.000 ;
    END
  END io_cpu_memory_mmuBus_cmd_virtualAddress[2]
  PIN io_cpu_memory_mmuBus_cmd_virtualAddress[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.930 246.000 577.210 250.000 ;
    END
  END io_cpu_memory_mmuBus_cmd_virtualAddress[30]
  PIN io_cpu_memory_mmuBus_cmd_virtualAddress[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.650 246.000 591.930 250.000 ;
    END
  END io_cpu_memory_mmuBus_cmd_virtualAddress[31]
  PIN io_cpu_memory_mmuBus_cmd_virtualAddress[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 246.000 165.050 250.000 ;
    END
  END io_cpu_memory_mmuBus_cmd_virtualAddress[3]
  PIN io_cpu_memory_mmuBus_cmd_virtualAddress[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.170 246.000 183.450 250.000 ;
    END
  END io_cpu_memory_mmuBus_cmd_virtualAddress[4]
  PIN io_cpu_memory_mmuBus_cmd_virtualAddress[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 246.000 200.010 250.000 ;
    END
  END io_cpu_memory_mmuBus_cmd_virtualAddress[5]
  PIN io_cpu_memory_mmuBus_cmd_virtualAddress[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 246.000 216.570 250.000 ;
    END
  END io_cpu_memory_mmuBus_cmd_virtualAddress[6]
  PIN io_cpu_memory_mmuBus_cmd_virtualAddress[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.850 246.000 233.130 250.000 ;
    END
  END io_cpu_memory_mmuBus_cmd_virtualAddress[7]
  PIN io_cpu_memory_mmuBus_cmd_virtualAddress[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 246.000 249.690 250.000 ;
    END
  END io_cpu_memory_mmuBus_cmd_virtualAddress[8]
  PIN io_cpu_memory_mmuBus_cmd_virtualAddress[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.970 246.000 266.250 250.000 ;
    END
  END io_cpu_memory_mmuBus_cmd_virtualAddress[9]
  PIN io_cpu_memory_mmuBus_end
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 246.000 69.370 250.000 ;
    END
  END io_cpu_memory_mmuBus_end
  PIN io_cpu_memory_mmuBus_rsp_allowExecute
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 246.000 71.210 250.000 ;
    END
  END io_cpu_memory_mmuBus_rsp_allowExecute
  PIN io_cpu_memory_mmuBus_rsp_allowRead
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 246.000 73.050 250.000 ;
    END
  END io_cpu_memory_mmuBus_rsp_allowRead
  PIN io_cpu_memory_mmuBus_rsp_allowWrite
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 246.000 74.890 250.000 ;
    END
  END io_cpu_memory_mmuBus_rsp_allowWrite
  PIN io_cpu_memory_mmuBus_rsp_exception
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 246.000 76.730 250.000 ;
    END
  END io_cpu_memory_mmuBus_rsp_exception
  PIN io_cpu_memory_mmuBus_rsp_isIoAccess
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 246.000 78.570 250.000 ;
    END
  END io_cpu_memory_mmuBus_rsp_isIoAccess
  PIN io_cpu_memory_mmuBus_rsp_physicalAddress[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 246.000 109.850 250.000 ;
    END
  END io_cpu_memory_mmuBus_rsp_physicalAddress[0]
  PIN io_cpu_memory_mmuBus_rsp_physicalAddress[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 246.000 284.650 250.000 ;
    END
  END io_cpu_memory_mmuBus_rsp_physicalAddress[10]
  PIN io_cpu_memory_mmuBus_rsp_physicalAddress[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.090 246.000 299.370 250.000 ;
    END
  END io_cpu_memory_mmuBus_rsp_physicalAddress[11]
  PIN io_cpu_memory_mmuBus_rsp_physicalAddress[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.810 246.000 314.090 250.000 ;
    END
  END io_cpu_memory_mmuBus_rsp_physicalAddress[12]
  PIN io_cpu_memory_mmuBus_rsp_physicalAddress[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 246.000 328.810 250.000 ;
    END
  END io_cpu_memory_mmuBus_rsp_physicalAddress[13]
  PIN io_cpu_memory_mmuBus_rsp_physicalAddress[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.250 246.000 343.530 250.000 ;
    END
  END io_cpu_memory_mmuBus_rsp_physicalAddress[14]
  PIN io_cpu_memory_mmuBus_rsp_physicalAddress[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.970 246.000 358.250 250.000 ;
    END
  END io_cpu_memory_mmuBus_rsp_physicalAddress[15]
  PIN io_cpu_memory_mmuBus_rsp_physicalAddress[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.690 246.000 372.970 250.000 ;
    END
  END io_cpu_memory_mmuBus_rsp_physicalAddress[16]
  PIN io_cpu_memory_mmuBus_rsp_physicalAddress[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.410 246.000 387.690 250.000 ;
    END
  END io_cpu_memory_mmuBus_rsp_physicalAddress[17]
  PIN io_cpu_memory_mmuBus_rsp_physicalAddress[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.130 246.000 402.410 250.000 ;
    END
  END io_cpu_memory_mmuBus_rsp_physicalAddress[18]
  PIN io_cpu_memory_mmuBus_rsp_physicalAddress[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.850 246.000 417.130 250.000 ;
    END
  END io_cpu_memory_mmuBus_rsp_physicalAddress[19]
  PIN io_cpu_memory_mmuBus_rsp_physicalAddress[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 246.000 130.090 250.000 ;
    END
  END io_cpu_memory_mmuBus_rsp_physicalAddress[1]
  PIN io_cpu_memory_mmuBus_rsp_physicalAddress[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 246.000 431.850 250.000 ;
    END
  END io_cpu_memory_mmuBus_rsp_physicalAddress[20]
  PIN io_cpu_memory_mmuBus_rsp_physicalAddress[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.290 246.000 446.570 250.000 ;
    END
  END io_cpu_memory_mmuBus_rsp_physicalAddress[21]
  PIN io_cpu_memory_mmuBus_rsp_physicalAddress[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.010 246.000 461.290 250.000 ;
    END
  END io_cpu_memory_mmuBus_rsp_physicalAddress[22]
  PIN io_cpu_memory_mmuBus_rsp_physicalAddress[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.730 246.000 476.010 250.000 ;
    END
  END io_cpu_memory_mmuBus_rsp_physicalAddress[23]
  PIN io_cpu_memory_mmuBus_rsp_physicalAddress[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.450 246.000 490.730 250.000 ;
    END
  END io_cpu_memory_mmuBus_rsp_physicalAddress[24]
  PIN io_cpu_memory_mmuBus_rsp_physicalAddress[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.170 246.000 505.450 250.000 ;
    END
  END io_cpu_memory_mmuBus_rsp_physicalAddress[25]
  PIN io_cpu_memory_mmuBus_rsp_physicalAddress[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.890 246.000 520.170 250.000 ;
    END
  END io_cpu_memory_mmuBus_rsp_physicalAddress[26]
  PIN io_cpu_memory_mmuBus_rsp_physicalAddress[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 246.000 534.890 250.000 ;
    END
  END io_cpu_memory_mmuBus_rsp_physicalAddress[27]
  PIN io_cpu_memory_mmuBus_rsp_physicalAddress[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.330 246.000 549.610 250.000 ;
    END
  END io_cpu_memory_mmuBus_rsp_physicalAddress[28]
  PIN io_cpu_memory_mmuBus_rsp_physicalAddress[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.050 246.000 564.330 250.000 ;
    END
  END io_cpu_memory_mmuBus_rsp_physicalAddress[29]
  PIN io_cpu_memory_mmuBus_rsp_physicalAddress[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 246.000 148.490 250.000 ;
    END
  END io_cpu_memory_mmuBus_rsp_physicalAddress[2]
  PIN io_cpu_memory_mmuBus_rsp_physicalAddress[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.770 246.000 579.050 250.000 ;
    END
  END io_cpu_memory_mmuBus_rsp_physicalAddress[30]
  PIN io_cpu_memory_mmuBus_rsp_physicalAddress[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.490 246.000 593.770 250.000 ;
    END
  END io_cpu_memory_mmuBus_rsp_physicalAddress[31]
  PIN io_cpu_memory_mmuBus_rsp_physicalAddress[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 246.000 166.890 250.000 ;
    END
  END io_cpu_memory_mmuBus_rsp_physicalAddress[3]
  PIN io_cpu_memory_mmuBus_rsp_physicalAddress[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 246.000 185.290 250.000 ;
    END
  END io_cpu_memory_mmuBus_rsp_physicalAddress[4]
  PIN io_cpu_memory_mmuBus_rsp_physicalAddress[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 246.000 201.850 250.000 ;
    END
  END io_cpu_memory_mmuBus_rsp_physicalAddress[5]
  PIN io_cpu_memory_mmuBus_rsp_physicalAddress[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 246.000 218.410 250.000 ;
    END
  END io_cpu_memory_mmuBus_rsp_physicalAddress[6]
  PIN io_cpu_memory_mmuBus_rsp_physicalAddress[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 246.000 234.970 250.000 ;
    END
  END io_cpu_memory_mmuBus_rsp_physicalAddress[7]
  PIN io_cpu_memory_mmuBus_rsp_physicalAddress[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 246.000 251.530 250.000 ;
    END
  END io_cpu_memory_mmuBus_rsp_physicalAddress[8]
  PIN io_cpu_memory_mmuBus_rsp_physicalAddress[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.810 246.000 268.090 250.000 ;
    END
  END io_cpu_memory_mmuBus_rsp_physicalAddress[9]
  PIN io_cpu_memory_mmuBus_rsp_refilling
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 246.000 80.410 250.000 ;
    END
  END io_cpu_memory_mmuBus_rsp_refilling
  PIN io_cpu_memory_mmuBus_spr_payload_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 246.000 111.690 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_payload_data[0]
  PIN io_cpu_memory_mmuBus_spr_payload_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.210 246.000 286.490 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_payload_data[10]
  PIN io_cpu_memory_mmuBus_spr_payload_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.930 246.000 301.210 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_payload_data[11]
  PIN io_cpu_memory_mmuBus_spr_payload_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 246.000 315.930 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_payload_data[12]
  PIN io_cpu_memory_mmuBus_spr_payload_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.370 246.000 330.650 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_payload_data[13]
  PIN io_cpu_memory_mmuBus_spr_payload_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 246.000 345.370 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_payload_data[14]
  PIN io_cpu_memory_mmuBus_spr_payload_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.810 246.000 360.090 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_payload_data[15]
  PIN io_cpu_memory_mmuBus_spr_payload_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 246.000 374.810 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_payload_data[16]
  PIN io_cpu_memory_mmuBus_spr_payload_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.250 246.000 389.530 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_payload_data[17]
  PIN io_cpu_memory_mmuBus_spr_payload_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.970 246.000 404.250 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_payload_data[18]
  PIN io_cpu_memory_mmuBus_spr_payload_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 246.000 418.970 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_payload_data[19]
  PIN io_cpu_memory_mmuBus_spr_payload_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 246.000 131.930 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_payload_data[1]
  PIN io_cpu_memory_mmuBus_spr_payload_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.410 246.000 433.690 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_payload_data[20]
  PIN io_cpu_memory_mmuBus_spr_payload_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.130 246.000 448.410 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_payload_data[21]
  PIN io_cpu_memory_mmuBus_spr_payload_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.850 246.000 463.130 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_payload_data[22]
  PIN io_cpu_memory_mmuBus_spr_payload_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.570 246.000 477.850 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_payload_data[23]
  PIN io_cpu_memory_mmuBus_spr_payload_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.290 246.000 492.570 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_payload_data[24]
  PIN io_cpu_memory_mmuBus_spr_payload_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.010 246.000 507.290 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_payload_data[25]
  PIN io_cpu_memory_mmuBus_spr_payload_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.730 246.000 522.010 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_payload_data[26]
  PIN io_cpu_memory_mmuBus_spr_payload_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.450 246.000 536.730 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_payload_data[27]
  PIN io_cpu_memory_mmuBus_spr_payload_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.170 246.000 551.450 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_payload_data[28]
  PIN io_cpu_memory_mmuBus_spr_payload_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.890 246.000 566.170 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_payload_data[29]
  PIN io_cpu_memory_mmuBus_spr_payload_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 246.000 150.330 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_payload_data[2]
  PIN io_cpu_memory_mmuBus_spr_payload_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.610 246.000 580.890 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_payload_data[30]
  PIN io_cpu_memory_mmuBus_spr_payload_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.330 246.000 595.610 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_payload_data[31]
  PIN io_cpu_memory_mmuBus_spr_payload_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 246.000 168.730 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_payload_data[3]
  PIN io_cpu_memory_mmuBus_spr_payload_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 246.000 187.130 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_payload_data[4]
  PIN io_cpu_memory_mmuBus_spr_payload_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 246.000 203.690 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_payload_data[5]
  PIN io_cpu_memory_mmuBus_spr_payload_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.970 246.000 220.250 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_payload_data[6]
  PIN io_cpu_memory_mmuBus_spr_payload_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.530 246.000 236.810 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_payload_data[7]
  PIN io_cpu_memory_mmuBus_spr_payload_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 246.000 253.370 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_payload_data[8]
  PIN io_cpu_memory_mmuBus_spr_payload_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 246.000 269.930 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_payload_data[9]
  PIN io_cpu_memory_mmuBus_spr_payload_id[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 246.000 113.530 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_payload_id[0]
  PIN io_cpu_memory_mmuBus_spr_payload_id[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 246.000 133.770 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_payload_id[1]
  PIN io_cpu_memory_mmuBus_spr_payload_id[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 246.000 152.170 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_payload_id[2]
  PIN io_cpu_memory_mmuBus_spr_payload_id[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 246.000 170.570 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_payload_id[3]
  PIN io_cpu_memory_mmuBus_spr_payload_id[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.690 246.000 188.970 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_payload_id[4]
  PIN io_cpu_memory_mmuBus_spr_payload_id[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 246.000 205.530 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_payload_id[5]
  PIN io_cpu_memory_mmuBus_spr_payload_id[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.810 246.000 222.090 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_payload_id[6]
  PIN io_cpu_memory_mmuBus_spr_payload_id[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 246.000 238.650 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_payload_id[7]
  PIN io_cpu_memory_mmuBus_spr_payload_id[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 246.000 255.210 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_payload_id[8]
  PIN io_cpu_memory_mmuBus_spr_payload_id[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.490 246.000 271.770 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_payload_id[9]
  PIN io_cpu_memory_mmuBus_spr_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 246.000 82.250 250.000 ;
    END
  END io_cpu_memory_mmuBus_spr_valid
  PIN io_cpu_redo
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 246.000 84.090 250.000 ;
    END
  END io_cpu_redo
  PIN io_cpu_writeBack_accessError
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 246.000 85.930 250.000 ;
    END
  END io_cpu_writeBack_accessError
  PIN io_cpu_writeBack_address[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 246.000 115.370 250.000 ;
    END
  END io_cpu_writeBack_address[0]
  PIN io_cpu_writeBack_address[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 246.000 288.330 250.000 ;
    END
  END io_cpu_writeBack_address[10]
  PIN io_cpu_writeBack_address[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 246.000 303.050 250.000 ;
    END
  END io_cpu_writeBack_address[11]
  PIN io_cpu_writeBack_address[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 246.000 317.770 250.000 ;
    END
  END io_cpu_writeBack_address[12]
  PIN io_cpu_writeBack_address[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.210 246.000 332.490 250.000 ;
    END
  END io_cpu_writeBack_address[13]
  PIN io_cpu_writeBack_address[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.930 246.000 347.210 250.000 ;
    END
  END io_cpu_writeBack_address[14]
  PIN io_cpu_writeBack_address[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.650 246.000 361.930 250.000 ;
    END
  END io_cpu_writeBack_address[15]
  PIN io_cpu_writeBack_address[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.370 246.000 376.650 250.000 ;
    END
  END io_cpu_writeBack_address[16]
  PIN io_cpu_writeBack_address[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.090 246.000 391.370 250.000 ;
    END
  END io_cpu_writeBack_address[17]
  PIN io_cpu_writeBack_address[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 246.000 406.090 250.000 ;
    END
  END io_cpu_writeBack_address[18]
  PIN io_cpu_writeBack_address[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.530 246.000 420.810 250.000 ;
    END
  END io_cpu_writeBack_address[19]
  PIN io_cpu_writeBack_address[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 246.000 135.610 250.000 ;
    END
  END io_cpu_writeBack_address[1]
  PIN io_cpu_writeBack_address[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.250 246.000 435.530 250.000 ;
    END
  END io_cpu_writeBack_address[20]
  PIN io_cpu_writeBack_address[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.970 246.000 450.250 250.000 ;
    END
  END io_cpu_writeBack_address[21]
  PIN io_cpu_writeBack_address[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.690 246.000 464.970 250.000 ;
    END
  END io_cpu_writeBack_address[22]
  PIN io_cpu_writeBack_address[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.410 246.000 479.690 250.000 ;
    END
  END io_cpu_writeBack_address[23]
  PIN io_cpu_writeBack_address[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.130 246.000 494.410 250.000 ;
    END
  END io_cpu_writeBack_address[24]
  PIN io_cpu_writeBack_address[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 246.000 509.130 250.000 ;
    END
  END io_cpu_writeBack_address[25]
  PIN io_cpu_writeBack_address[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.570 246.000 523.850 250.000 ;
    END
  END io_cpu_writeBack_address[26]
  PIN io_cpu_writeBack_address[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.290 246.000 538.570 250.000 ;
    END
  END io_cpu_writeBack_address[27]
  PIN io_cpu_writeBack_address[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.010 246.000 553.290 250.000 ;
    END
  END io_cpu_writeBack_address[28]
  PIN io_cpu_writeBack_address[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.730 246.000 568.010 250.000 ;
    END
  END io_cpu_writeBack_address[29]
  PIN io_cpu_writeBack_address[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 246.000 154.010 250.000 ;
    END
  END io_cpu_writeBack_address[2]
  PIN io_cpu_writeBack_address[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.450 246.000 582.730 250.000 ;
    END
  END io_cpu_writeBack_address[30]
  PIN io_cpu_writeBack_address[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.170 246.000 597.450 250.000 ;
    END
  END io_cpu_writeBack_address[31]
  PIN io_cpu_writeBack_address[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.130 246.000 172.410 250.000 ;
    END
  END io_cpu_writeBack_address[3]
  PIN io_cpu_writeBack_address[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 246.000 190.810 250.000 ;
    END
  END io_cpu_writeBack_address[4]
  PIN io_cpu_writeBack_address[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 246.000 207.370 250.000 ;
    END
  END io_cpu_writeBack_address[5]
  PIN io_cpu_writeBack_address[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.650 246.000 223.930 250.000 ;
    END
  END io_cpu_writeBack_address[6]
  PIN io_cpu_writeBack_address[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 246.000 240.490 250.000 ;
    END
  END io_cpu_writeBack_address[7]
  PIN io_cpu_writeBack_address[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.770 246.000 257.050 250.000 ;
    END
  END io_cpu_writeBack_address[8]
  PIN io_cpu_writeBack_address[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 246.000 273.610 250.000 ;
    END
  END io_cpu_writeBack_address[9]
  PIN io_cpu_writeBack_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 246.000 117.210 250.000 ;
    END
  END io_cpu_writeBack_data[0]
  PIN io_cpu_writeBack_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 246.000 290.170 250.000 ;
    END
  END io_cpu_writeBack_data[10]
  PIN io_cpu_writeBack_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.610 246.000 304.890 250.000 ;
    END
  END io_cpu_writeBack_data[11]
  PIN io_cpu_writeBack_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 246.000 319.610 250.000 ;
    END
  END io_cpu_writeBack_data[12]
  PIN io_cpu_writeBack_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 246.000 334.330 250.000 ;
    END
  END io_cpu_writeBack_data[13]
  PIN io_cpu_writeBack_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.770 246.000 349.050 250.000 ;
    END
  END io_cpu_writeBack_data[14]
  PIN io_cpu_writeBack_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 246.000 363.770 250.000 ;
    END
  END io_cpu_writeBack_data[15]
  PIN io_cpu_writeBack_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 246.000 378.490 250.000 ;
    END
  END io_cpu_writeBack_data[16]
  PIN io_cpu_writeBack_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 246.000 393.210 250.000 ;
    END
  END io_cpu_writeBack_data[17]
  PIN io_cpu_writeBack_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.650 246.000 407.930 250.000 ;
    END
  END io_cpu_writeBack_data[18]
  PIN io_cpu_writeBack_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.370 246.000 422.650 250.000 ;
    END
  END io_cpu_writeBack_data[19]
  PIN io_cpu_writeBack_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 246.000 137.450 250.000 ;
    END
  END io_cpu_writeBack_data[1]
  PIN io_cpu_writeBack_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.090 246.000 437.370 250.000 ;
    END
  END io_cpu_writeBack_data[20]
  PIN io_cpu_writeBack_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.810 246.000 452.090 250.000 ;
    END
  END io_cpu_writeBack_data[21]
  PIN io_cpu_writeBack_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.530 246.000 466.810 250.000 ;
    END
  END io_cpu_writeBack_data[22]
  PIN io_cpu_writeBack_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.250 246.000 481.530 250.000 ;
    END
  END io_cpu_writeBack_data[23]
  PIN io_cpu_writeBack_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 246.000 496.250 250.000 ;
    END
  END io_cpu_writeBack_data[24]
  PIN io_cpu_writeBack_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.690 246.000 510.970 250.000 ;
    END
  END io_cpu_writeBack_data[25]
  PIN io_cpu_writeBack_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.410 246.000 525.690 250.000 ;
    END
  END io_cpu_writeBack_data[26]
  PIN io_cpu_writeBack_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.130 246.000 540.410 250.000 ;
    END
  END io_cpu_writeBack_data[27]
  PIN io_cpu_writeBack_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.850 246.000 555.130 250.000 ;
    END
  END io_cpu_writeBack_data[28]
  PIN io_cpu_writeBack_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.570 246.000 569.850 250.000 ;
    END
  END io_cpu_writeBack_data[29]
  PIN io_cpu_writeBack_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 246.000 155.850 250.000 ;
    END
  END io_cpu_writeBack_data[2]
  PIN io_cpu_writeBack_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.290 246.000 584.570 250.000 ;
    END
  END io_cpu_writeBack_data[30]
  PIN io_cpu_writeBack_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 246.000 599.290 250.000 ;
    END
  END io_cpu_writeBack_data[31]
  PIN io_cpu_writeBack_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 246.000 174.250 250.000 ;
    END
  END io_cpu_writeBack_data[3]
  PIN io_cpu_writeBack_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 246.000 192.650 250.000 ;
    END
  END io_cpu_writeBack_data[4]
  PIN io_cpu_writeBack_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 246.000 209.210 250.000 ;
    END
  END io_cpu_writeBack_data[5]
  PIN io_cpu_writeBack_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 246.000 225.770 250.000 ;
    END
  END io_cpu_writeBack_data[6]
  PIN io_cpu_writeBack_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 246.000 242.330 250.000 ;
    END
  END io_cpu_writeBack_data[7]
  PIN io_cpu_writeBack_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 246.000 258.890 250.000 ;
    END
  END io_cpu_writeBack_data[8]
  PIN io_cpu_writeBack_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.170 246.000 275.450 250.000 ;
    END
  END io_cpu_writeBack_data[9]
  PIN io_cpu_writeBack_exceptionType[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 246.000 119.050 250.000 ;
    END
  END io_cpu_writeBack_exceptionType[0]
  PIN io_cpu_writeBack_exceptionType[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 246.000 139.290 250.000 ;
    END
  END io_cpu_writeBack_exceptionType[1]
  PIN io_cpu_writeBack_exceptionType[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 246.000 157.690 250.000 ;
    END
  END io_cpu_writeBack_exceptionType[2]
  PIN io_cpu_writeBack_exceptionType[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 246.000 176.090 250.000 ;
    END
  END io_cpu_writeBack_exceptionType[3]
  PIN io_cpu_writeBack_haltIt
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 246.000 87.770 250.000 ;
    END
  END io_cpu_writeBack_haltIt
  PIN io_cpu_writeBack_isStuck
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 246.000 89.610 250.000 ;
    END
  END io_cpu_writeBack_isStuck
  PIN io_cpu_writeBack_isUser
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 246.000 91.450 250.000 ;
    END
  END io_cpu_writeBack_isUser
  PIN io_cpu_writeBack_isValid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 246.000 93.290 250.000 ;
    END
  END io_cpu_writeBack_isValid
  PIN io_cpu_writeBack_isWrite
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 246.000 95.130 250.000 ;
    END
  END io_cpu_writeBack_isWrite
  PIN io_cpu_writeBack_mmuException
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 246.000 96.970 250.000 ;
    END
  END io_cpu_writeBack_mmuException
  PIN io_cpu_writeBack_unalignedAccess
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 246.000 98.810 250.000 ;
    END
  END io_cpu_writeBack_unalignedAccess
  PIN io_mem_cmd_payload_address[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END io_mem_cmd_payload_address[0]
  PIN io_mem_cmd_payload_address[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END io_mem_cmd_payload_address[10]
  PIN io_mem_cmd_payload_address[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 0.000 280.970 4.000 ;
    END
  END io_mem_cmd_payload_address[11]
  PIN io_mem_cmd_payload_address[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 0.000 297.530 4.000 ;
    END
  END io_mem_cmd_payload_address[12]
  PIN io_mem_cmd_payload_address[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.810 0.000 314.090 4.000 ;
    END
  END io_mem_cmd_payload_address[13]
  PIN io_mem_cmd_payload_address[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.370 0.000 330.650 4.000 ;
    END
  END io_mem_cmd_payload_address[14]
  PIN io_mem_cmd_payload_address[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.930 0.000 347.210 4.000 ;
    END
  END io_mem_cmd_payload_address[15]
  PIN io_mem_cmd_payload_address[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 0.000 363.770 4.000 ;
    END
  END io_mem_cmd_payload_address[16]
  PIN io_mem_cmd_payload_address[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 0.000 380.330 4.000 ;
    END
  END io_mem_cmd_payload_address[17]
  PIN io_mem_cmd_payload_address[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.610 0.000 396.890 4.000 ;
    END
  END io_mem_cmd_payload_address[18]
  PIN io_mem_cmd_payload_address[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.170 0.000 413.450 4.000 ;
    END
  END io_mem_cmd_payload_address[19]
  PIN io_mem_cmd_payload_address[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END io_mem_cmd_payload_address[1]
  PIN io_mem_cmd_payload_address[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.730 0.000 430.010 4.000 ;
    END
  END io_mem_cmd_payload_address[20]
  PIN io_mem_cmd_payload_address[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.290 0.000 446.570 4.000 ;
    END
  END io_mem_cmd_payload_address[21]
  PIN io_mem_cmd_payload_address[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.850 0.000 463.130 4.000 ;
    END
  END io_mem_cmd_payload_address[22]
  PIN io_mem_cmd_payload_address[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.410 0.000 479.690 4.000 ;
    END
  END io_mem_cmd_payload_address[23]
  PIN io_mem_cmd_payload_address[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 0.000 496.250 4.000 ;
    END
  END io_mem_cmd_payload_address[24]
  PIN io_mem_cmd_payload_address[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.530 0.000 512.810 4.000 ;
    END
  END io_mem_cmd_payload_address[25]
  PIN io_mem_cmd_payload_address[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.090 0.000 529.370 4.000 ;
    END
  END io_mem_cmd_payload_address[26]
  PIN io_mem_cmd_payload_address[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.650 0.000 545.930 4.000 ;
    END
  END io_mem_cmd_payload_address[27]
  PIN io_mem_cmd_payload_address[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.210 0.000 562.490 4.000 ;
    END
  END io_mem_cmd_payload_address[28]
  PIN io_mem_cmd_payload_address[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.770 0.000 579.050 4.000 ;
    END
  END io_mem_cmd_payload_address[29]
  PIN io_mem_cmd_payload_address[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END io_mem_cmd_payload_address[2]
  PIN io_mem_cmd_payload_address[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.330 0.000 595.610 4.000 ;
    END
  END io_mem_cmd_payload_address[30]
  PIN io_mem_cmd_payload_address[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.890 0.000 612.170 4.000 ;
    END
  END io_mem_cmd_payload_address[31]
  PIN io_mem_cmd_payload_address[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END io_mem_cmd_payload_address[3]
  PIN io_mem_cmd_payload_address[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 0.000 165.050 4.000 ;
    END
  END io_mem_cmd_payload_address[4]
  PIN io_mem_cmd_payload_address[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.330 0.000 181.610 4.000 ;
    END
  END io_mem_cmd_payload_address[5]
  PIN io_mem_cmd_payload_address[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 0.000 198.170 4.000 ;
    END
  END io_mem_cmd_payload_address[6]
  PIN io_mem_cmd_payload_address[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 0.000 214.730 4.000 ;
    END
  END io_mem_cmd_payload_address[7]
  PIN io_mem_cmd_payload_address[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 4.000 ;
    END
  END io_mem_cmd_payload_address[8]
  PIN io_mem_cmd_payload_address[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.570 0.000 247.850 4.000 ;
    END
  END io_mem_cmd_payload_address[9]
  PIN io_mem_cmd_payload_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 4.000 ;
    END
  END io_mem_cmd_payload_data[0]
  PIN io_mem_cmd_payload_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 0.000 269.930 4.000 ;
    END
  END io_mem_cmd_payload_data[10]
  PIN io_mem_cmd_payload_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.210 0.000 286.490 4.000 ;
    END
  END io_mem_cmd_payload_data[11]
  PIN io_mem_cmd_payload_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END io_mem_cmd_payload_data[12]
  PIN io_mem_cmd_payload_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 0.000 319.610 4.000 ;
    END
  END io_mem_cmd_payload_data[13]
  PIN io_mem_cmd_payload_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.890 0.000 336.170 4.000 ;
    END
  END io_mem_cmd_payload_data[14]
  PIN io_mem_cmd_payload_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.450 0.000 352.730 4.000 ;
    END
  END io_mem_cmd_payload_data[15]
  PIN io_mem_cmd_payload_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.010 0.000 369.290 4.000 ;
    END
  END io_mem_cmd_payload_data[16]
  PIN io_mem_cmd_payload_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.570 0.000 385.850 4.000 ;
    END
  END io_mem_cmd_payload_data[17]
  PIN io_mem_cmd_payload_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.130 0.000 402.410 4.000 ;
    END
  END io_mem_cmd_payload_data[18]
  PIN io_mem_cmd_payload_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 0.000 418.970 4.000 ;
    END
  END io_mem_cmd_payload_data[19]
  PIN io_mem_cmd_payload_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END io_mem_cmd_payload_data[1]
  PIN io_mem_cmd_payload_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.250 0.000 435.530 4.000 ;
    END
  END io_mem_cmd_payload_data[20]
  PIN io_mem_cmd_payload_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.810 0.000 452.090 4.000 ;
    END
  END io_mem_cmd_payload_data[21]
  PIN io_mem_cmd_payload_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.370 0.000 468.650 4.000 ;
    END
  END io_mem_cmd_payload_data[22]
  PIN io_mem_cmd_payload_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.930 0.000 485.210 4.000 ;
    END
  END io_mem_cmd_payload_data[23]
  PIN io_mem_cmd_payload_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.490 0.000 501.770 4.000 ;
    END
  END io_mem_cmd_payload_data[24]
  PIN io_mem_cmd_payload_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.050 0.000 518.330 4.000 ;
    END
  END io_mem_cmd_payload_data[25]
  PIN io_mem_cmd_payload_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 0.000 534.890 4.000 ;
    END
  END io_mem_cmd_payload_data[26]
  PIN io_mem_cmd_payload_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.170 0.000 551.450 4.000 ;
    END
  END io_mem_cmd_payload_data[27]
  PIN io_mem_cmd_payload_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.730 0.000 568.010 4.000 ;
    END
  END io_mem_cmd_payload_data[28]
  PIN io_mem_cmd_payload_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.290 0.000 584.570 4.000 ;
    END
  END io_mem_cmd_payload_data[29]
  PIN io_mem_cmd_payload_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END io_mem_cmd_payload_data[2]
  PIN io_mem_cmd_payload_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 600.850 0.000 601.130 4.000 ;
    END
  END io_mem_cmd_payload_data[30]
  PIN io_mem_cmd_payload_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.410 0.000 617.690 4.000 ;
    END
  END io_mem_cmd_payload_data[31]
  PIN io_mem_cmd_payload_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END io_mem_cmd_payload_data[3]
  PIN io_mem_cmd_payload_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 4.000 ;
    END
  END io_mem_cmd_payload_data[4]
  PIN io_mem_cmd_payload_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END io_mem_cmd_payload_data[5]
  PIN io_mem_cmd_payload_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 0.000 203.690 4.000 ;
    END
  END io_mem_cmd_payload_data[6]
  PIN io_mem_cmd_payload_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.970 0.000 220.250 4.000 ;
    END
  END io_mem_cmd_payload_data[7]
  PIN io_mem_cmd_payload_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.530 0.000 236.810 4.000 ;
    END
  END io_mem_cmd_payload_data[8]
  PIN io_mem_cmd_payload_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 0.000 253.370 4.000 ;
    END
  END io_mem_cmd_payload_data[9]
  PIN io_mem_cmd_payload_last
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 4.000 ;
    END
  END io_mem_cmd_payload_last
  PIN io_mem_cmd_payload_length[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END io_mem_cmd_payload_length[0]
  PIN io_mem_cmd_payload_length[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 4.000 ;
    END
  END io_mem_cmd_payload_length[1]
  PIN io_mem_cmd_payload_length[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 4.000 ;
    END
  END io_mem_cmd_payload_length[2]
  PIN io_mem_cmd_payload_mask[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 4.000 ;
    END
  END io_mem_cmd_payload_mask[0]
  PIN io_mem_cmd_payload_mask[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 4.000 ;
    END
  END io_mem_cmd_payload_mask[1]
  PIN io_mem_cmd_payload_mask[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 0.000 131.930 4.000 ;
    END
  END io_mem_cmd_payload_mask[2]
  PIN io_mem_cmd_payload_mask[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 0.000 154.010 4.000 ;
    END
  END io_mem_cmd_payload_mask[3]
  PIN io_mem_cmd_payload_wr
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END io_mem_cmd_payload_wr
  PIN io_mem_cmd_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 4.000 ;
    END
  END io_mem_cmd_ready
  PIN io_mem_cmd_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END io_mem_cmd_valid
  PIN io_mem_rsp_payload_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 4.000 ;
    END
  END io_mem_rsp_payload_data[0]
  PIN io_mem_rsp_payload_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.170 0.000 275.450 4.000 ;
    END
  END io_mem_rsp_payload_data[10]
  PIN io_mem_rsp_payload_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.730 0.000 292.010 4.000 ;
    END
  END io_mem_rsp_payload_data[11]
  PIN io_mem_rsp_payload_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 0.000 308.570 4.000 ;
    END
  END io_mem_rsp_payload_data[12]
  PIN io_mem_rsp_payload_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.850 0.000 325.130 4.000 ;
    END
  END io_mem_rsp_payload_data[13]
  PIN io_mem_rsp_payload_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END io_mem_rsp_payload_data[14]
  PIN io_mem_rsp_payload_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.970 0.000 358.250 4.000 ;
    END
  END io_mem_rsp_payload_data[15]
  PIN io_mem_rsp_payload_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 0.000 374.810 4.000 ;
    END
  END io_mem_rsp_payload_data[16]
  PIN io_mem_rsp_payload_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.090 0.000 391.370 4.000 ;
    END
  END io_mem_rsp_payload_data[17]
  PIN io_mem_rsp_payload_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.650 0.000 407.930 4.000 ;
    END
  END io_mem_rsp_payload_data[18]
  PIN io_mem_rsp_payload_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.210 0.000 424.490 4.000 ;
    END
  END io_mem_rsp_payload_data[19]
  PIN io_mem_rsp_payload_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END io_mem_rsp_payload_data[1]
  PIN io_mem_rsp_payload_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.770 0.000 441.050 4.000 ;
    END
  END io_mem_rsp_payload_data[20]
  PIN io_mem_rsp_payload_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 0.000 457.610 4.000 ;
    END
  END io_mem_rsp_payload_data[21]
  PIN io_mem_rsp_payload_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.890 0.000 474.170 4.000 ;
    END
  END io_mem_rsp_payload_data[22]
  PIN io_mem_rsp_payload_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.450 0.000 490.730 4.000 ;
    END
  END io_mem_rsp_payload_data[23]
  PIN io_mem_rsp_payload_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.010 0.000 507.290 4.000 ;
    END
  END io_mem_rsp_payload_data[24]
  PIN io_mem_rsp_payload_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.570 0.000 523.850 4.000 ;
    END
  END io_mem_rsp_payload_data[25]
  PIN io_mem_rsp_payload_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.130 0.000 540.410 4.000 ;
    END
  END io_mem_rsp_payload_data[26]
  PIN io_mem_rsp_payload_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 0.000 556.970 4.000 ;
    END
  END io_mem_rsp_payload_data[27]
  PIN io_mem_rsp_payload_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 0.000 573.530 4.000 ;
    END
  END io_mem_rsp_payload_data[28]
  PIN io_mem_rsp_payload_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.810 0.000 590.090 4.000 ;
    END
  END io_mem_rsp_payload_data[29]
  PIN io_mem_rsp_payload_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 4.000 ;
    END
  END io_mem_rsp_payload_data[2]
  PIN io_mem_rsp_payload_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.370 0.000 606.650 4.000 ;
    END
  END io_mem_rsp_payload_data[30]
  PIN io_mem_rsp_payload_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.930 0.000 623.210 4.000 ;
    END
  END io_mem_rsp_payload_data[31]
  PIN io_mem_rsp_payload_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 0.000 159.530 4.000 ;
    END
  END io_mem_rsp_payload_data[3]
  PIN io_mem_rsp_payload_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 0.000 176.090 4.000 ;
    END
  END io_mem_rsp_payload_data[4]
  PIN io_mem_rsp_payload_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 4.000 ;
    END
  END io_mem_rsp_payload_data[5]
  PIN io_mem_rsp_payload_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 0.000 209.210 4.000 ;
    END
  END io_mem_rsp_payload_data[6]
  PIN io_mem_rsp_payload_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END io_mem_rsp_payload_data[7]
  PIN io_mem_rsp_payload_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 0.000 242.330 4.000 ;
    END
  END io_mem_rsp_payload_data[8]
  PIN io_mem_rsp_payload_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 4.000 ;
    END
  END io_mem_rsp_payload_data[9]
  PIN io_mem_rsp_payload_error
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END io_mem_rsp_payload_error
  PIN io_mem_rsp_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 0.000 54.650 4.000 ;
    END
  END io_mem_rsp_valid
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.690 246.000 602.970 250.000 ;
    END
  END reset
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 179.160 22.640 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 179.160 176.240 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 179.160 329.840 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 179.160 483.440 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 7.940 10.640 9.540 182.480 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 179.160 99.440 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 179.160 253.040 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 179.160 406.640 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 179.160 560.240 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 10.700 10.640 12.300 182.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 630.780 10.640 632.380 179.760 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 644.460 236.725 ;
      LAYER met1 ;
        RECT 0.070 0.040 644.460 247.820 ;
      LAYER met2 ;
        RECT 0.100 245.720 46.730 247.850 ;
        RECT 47.570 245.720 48.570 247.850 ;
        RECT 49.410 245.720 50.410 247.850 ;
        RECT 51.250 245.720 52.250 247.850 ;
        RECT 53.090 245.720 54.090 247.850 ;
        RECT 54.930 245.720 55.930 247.850 ;
        RECT 56.770 245.720 57.770 247.850 ;
        RECT 58.610 245.720 59.610 247.850 ;
        RECT 60.450 245.720 61.450 247.850 ;
        RECT 62.290 245.720 63.290 247.850 ;
        RECT 64.130 245.720 65.130 247.850 ;
        RECT 65.970 245.720 66.970 247.850 ;
        RECT 67.810 245.720 68.810 247.850 ;
        RECT 69.650 245.720 70.650 247.850 ;
        RECT 71.490 245.720 72.490 247.850 ;
        RECT 73.330 245.720 74.330 247.850 ;
        RECT 75.170 245.720 76.170 247.850 ;
        RECT 77.010 245.720 78.010 247.850 ;
        RECT 78.850 245.720 79.850 247.850 ;
        RECT 80.690 245.720 81.690 247.850 ;
        RECT 82.530 245.720 83.530 247.850 ;
        RECT 84.370 245.720 85.370 247.850 ;
        RECT 86.210 245.720 87.210 247.850 ;
        RECT 88.050 245.720 89.050 247.850 ;
        RECT 89.890 245.720 90.890 247.850 ;
        RECT 91.730 245.720 92.730 247.850 ;
        RECT 93.570 245.720 94.570 247.850 ;
        RECT 95.410 245.720 96.410 247.850 ;
        RECT 97.250 245.720 98.250 247.850 ;
        RECT 99.090 245.720 100.090 247.850 ;
        RECT 100.930 245.720 101.930 247.850 ;
        RECT 102.770 245.720 103.770 247.850 ;
        RECT 104.610 245.720 105.610 247.850 ;
        RECT 106.450 245.720 107.450 247.850 ;
        RECT 108.290 245.720 109.290 247.850 ;
        RECT 110.130 245.720 111.130 247.850 ;
        RECT 111.970 245.720 112.970 247.850 ;
        RECT 113.810 245.720 114.810 247.850 ;
        RECT 115.650 245.720 116.650 247.850 ;
        RECT 117.490 245.720 118.490 247.850 ;
        RECT 119.330 245.720 120.330 247.850 ;
        RECT 121.170 245.720 122.170 247.850 ;
        RECT 123.010 245.720 124.010 247.850 ;
        RECT 124.850 245.720 125.850 247.850 ;
        RECT 126.690 245.720 127.690 247.850 ;
        RECT 128.530 245.720 129.530 247.850 ;
        RECT 130.370 245.720 131.370 247.850 ;
        RECT 132.210 245.720 133.210 247.850 ;
        RECT 134.050 245.720 135.050 247.850 ;
        RECT 135.890 245.720 136.890 247.850 ;
        RECT 137.730 245.720 138.730 247.850 ;
        RECT 139.570 245.720 140.570 247.850 ;
        RECT 141.410 245.720 142.410 247.850 ;
        RECT 143.250 245.720 144.250 247.850 ;
        RECT 145.090 245.720 146.090 247.850 ;
        RECT 146.930 245.720 147.930 247.850 ;
        RECT 148.770 245.720 149.770 247.850 ;
        RECT 150.610 245.720 151.610 247.850 ;
        RECT 152.450 245.720 153.450 247.850 ;
        RECT 154.290 245.720 155.290 247.850 ;
        RECT 156.130 245.720 157.130 247.850 ;
        RECT 157.970 245.720 158.970 247.850 ;
        RECT 159.810 245.720 160.810 247.850 ;
        RECT 161.650 245.720 162.650 247.850 ;
        RECT 163.490 245.720 164.490 247.850 ;
        RECT 165.330 245.720 166.330 247.850 ;
        RECT 167.170 245.720 168.170 247.850 ;
        RECT 169.010 245.720 170.010 247.850 ;
        RECT 170.850 245.720 171.850 247.850 ;
        RECT 172.690 245.720 173.690 247.850 ;
        RECT 174.530 245.720 175.530 247.850 ;
        RECT 176.370 245.720 177.370 247.850 ;
        RECT 178.210 245.720 179.210 247.850 ;
        RECT 180.050 245.720 181.050 247.850 ;
        RECT 181.890 245.720 182.890 247.850 ;
        RECT 183.730 245.720 184.730 247.850 ;
        RECT 185.570 245.720 186.570 247.850 ;
        RECT 187.410 245.720 188.410 247.850 ;
        RECT 189.250 245.720 190.250 247.850 ;
        RECT 191.090 245.720 192.090 247.850 ;
        RECT 192.930 245.720 193.930 247.850 ;
        RECT 194.770 245.720 195.770 247.850 ;
        RECT 196.610 245.720 197.610 247.850 ;
        RECT 198.450 245.720 199.450 247.850 ;
        RECT 200.290 245.720 201.290 247.850 ;
        RECT 202.130 245.720 203.130 247.850 ;
        RECT 203.970 245.720 204.970 247.850 ;
        RECT 205.810 245.720 206.810 247.850 ;
        RECT 207.650 245.720 208.650 247.850 ;
        RECT 209.490 245.720 210.490 247.850 ;
        RECT 211.330 245.720 212.330 247.850 ;
        RECT 213.170 245.720 214.170 247.850 ;
        RECT 215.010 245.720 216.010 247.850 ;
        RECT 216.850 245.720 217.850 247.850 ;
        RECT 218.690 245.720 219.690 247.850 ;
        RECT 220.530 245.720 221.530 247.850 ;
        RECT 222.370 245.720 223.370 247.850 ;
        RECT 224.210 245.720 225.210 247.850 ;
        RECT 226.050 245.720 227.050 247.850 ;
        RECT 227.890 245.720 228.890 247.850 ;
        RECT 229.730 245.720 230.730 247.850 ;
        RECT 231.570 245.720 232.570 247.850 ;
        RECT 233.410 245.720 234.410 247.850 ;
        RECT 235.250 245.720 236.250 247.850 ;
        RECT 237.090 245.720 238.090 247.850 ;
        RECT 238.930 245.720 239.930 247.850 ;
        RECT 240.770 245.720 241.770 247.850 ;
        RECT 242.610 245.720 243.610 247.850 ;
        RECT 244.450 245.720 245.450 247.850 ;
        RECT 246.290 245.720 247.290 247.850 ;
        RECT 248.130 245.720 249.130 247.850 ;
        RECT 249.970 245.720 250.970 247.850 ;
        RECT 251.810 245.720 252.810 247.850 ;
        RECT 253.650 245.720 254.650 247.850 ;
        RECT 255.490 245.720 256.490 247.850 ;
        RECT 257.330 245.720 258.330 247.850 ;
        RECT 259.170 245.720 260.170 247.850 ;
        RECT 261.010 245.720 262.010 247.850 ;
        RECT 262.850 245.720 263.850 247.850 ;
        RECT 264.690 245.720 265.690 247.850 ;
        RECT 266.530 245.720 267.530 247.850 ;
        RECT 268.370 245.720 269.370 247.850 ;
        RECT 270.210 245.720 271.210 247.850 ;
        RECT 272.050 245.720 273.050 247.850 ;
        RECT 273.890 245.720 274.890 247.850 ;
        RECT 275.730 245.720 276.730 247.850 ;
        RECT 277.570 245.720 278.570 247.850 ;
        RECT 279.410 245.720 280.410 247.850 ;
        RECT 281.250 245.720 282.250 247.850 ;
        RECT 283.090 245.720 284.090 247.850 ;
        RECT 284.930 245.720 285.930 247.850 ;
        RECT 286.770 245.720 287.770 247.850 ;
        RECT 288.610 245.720 289.610 247.850 ;
        RECT 290.450 245.720 291.450 247.850 ;
        RECT 292.290 245.720 293.290 247.850 ;
        RECT 294.130 245.720 295.130 247.850 ;
        RECT 295.970 245.720 296.970 247.850 ;
        RECT 297.810 245.720 298.810 247.850 ;
        RECT 299.650 245.720 300.650 247.850 ;
        RECT 301.490 245.720 302.490 247.850 ;
        RECT 303.330 245.720 304.330 247.850 ;
        RECT 305.170 245.720 306.170 247.850 ;
        RECT 307.010 245.720 308.010 247.850 ;
        RECT 308.850 245.720 309.850 247.850 ;
        RECT 310.690 245.720 311.690 247.850 ;
        RECT 312.530 245.720 313.530 247.850 ;
        RECT 314.370 245.720 315.370 247.850 ;
        RECT 316.210 245.720 317.210 247.850 ;
        RECT 318.050 245.720 319.050 247.850 ;
        RECT 319.890 245.720 320.890 247.850 ;
        RECT 321.730 245.720 322.730 247.850 ;
        RECT 323.570 245.720 324.570 247.850 ;
        RECT 325.410 245.720 326.410 247.850 ;
        RECT 327.250 245.720 328.250 247.850 ;
        RECT 329.090 245.720 330.090 247.850 ;
        RECT 330.930 245.720 331.930 247.850 ;
        RECT 332.770 245.720 333.770 247.850 ;
        RECT 334.610 245.720 335.610 247.850 ;
        RECT 336.450 245.720 337.450 247.850 ;
        RECT 338.290 245.720 339.290 247.850 ;
        RECT 340.130 245.720 341.130 247.850 ;
        RECT 341.970 245.720 342.970 247.850 ;
        RECT 343.810 245.720 344.810 247.850 ;
        RECT 345.650 245.720 346.650 247.850 ;
        RECT 347.490 245.720 348.490 247.850 ;
        RECT 349.330 245.720 350.330 247.850 ;
        RECT 351.170 245.720 352.170 247.850 ;
        RECT 353.010 245.720 354.010 247.850 ;
        RECT 354.850 245.720 355.850 247.850 ;
        RECT 356.690 245.720 357.690 247.850 ;
        RECT 358.530 245.720 359.530 247.850 ;
        RECT 360.370 245.720 361.370 247.850 ;
        RECT 362.210 245.720 363.210 247.850 ;
        RECT 364.050 245.720 365.050 247.850 ;
        RECT 365.890 245.720 366.890 247.850 ;
        RECT 367.730 245.720 368.730 247.850 ;
        RECT 369.570 245.720 370.570 247.850 ;
        RECT 371.410 245.720 372.410 247.850 ;
        RECT 373.250 245.720 374.250 247.850 ;
        RECT 375.090 245.720 376.090 247.850 ;
        RECT 376.930 245.720 377.930 247.850 ;
        RECT 378.770 245.720 379.770 247.850 ;
        RECT 380.610 245.720 381.610 247.850 ;
        RECT 382.450 245.720 383.450 247.850 ;
        RECT 384.290 245.720 385.290 247.850 ;
        RECT 386.130 245.720 387.130 247.850 ;
        RECT 387.970 245.720 388.970 247.850 ;
        RECT 389.810 245.720 390.810 247.850 ;
        RECT 391.650 245.720 392.650 247.850 ;
        RECT 393.490 245.720 394.490 247.850 ;
        RECT 395.330 245.720 396.330 247.850 ;
        RECT 397.170 245.720 398.170 247.850 ;
        RECT 399.010 245.720 400.010 247.850 ;
        RECT 400.850 245.720 401.850 247.850 ;
        RECT 402.690 245.720 403.690 247.850 ;
        RECT 404.530 245.720 405.530 247.850 ;
        RECT 406.370 245.720 407.370 247.850 ;
        RECT 408.210 245.720 409.210 247.850 ;
        RECT 410.050 245.720 411.050 247.850 ;
        RECT 411.890 245.720 412.890 247.850 ;
        RECT 413.730 245.720 414.730 247.850 ;
        RECT 415.570 245.720 416.570 247.850 ;
        RECT 417.410 245.720 418.410 247.850 ;
        RECT 419.250 245.720 420.250 247.850 ;
        RECT 421.090 245.720 422.090 247.850 ;
        RECT 422.930 245.720 423.930 247.850 ;
        RECT 424.770 245.720 425.770 247.850 ;
        RECT 426.610 245.720 427.610 247.850 ;
        RECT 428.450 245.720 429.450 247.850 ;
        RECT 430.290 245.720 431.290 247.850 ;
        RECT 432.130 245.720 433.130 247.850 ;
        RECT 433.970 245.720 434.970 247.850 ;
        RECT 435.810 245.720 436.810 247.850 ;
        RECT 437.650 245.720 438.650 247.850 ;
        RECT 439.490 245.720 440.490 247.850 ;
        RECT 441.330 245.720 442.330 247.850 ;
        RECT 443.170 245.720 444.170 247.850 ;
        RECT 445.010 245.720 446.010 247.850 ;
        RECT 446.850 245.720 447.850 247.850 ;
        RECT 448.690 245.720 449.690 247.850 ;
        RECT 450.530 245.720 451.530 247.850 ;
        RECT 452.370 245.720 453.370 247.850 ;
        RECT 454.210 245.720 455.210 247.850 ;
        RECT 456.050 245.720 457.050 247.850 ;
        RECT 457.890 245.720 458.890 247.850 ;
        RECT 459.730 245.720 460.730 247.850 ;
        RECT 461.570 245.720 462.570 247.850 ;
        RECT 463.410 245.720 464.410 247.850 ;
        RECT 465.250 245.720 466.250 247.850 ;
        RECT 467.090 245.720 468.090 247.850 ;
        RECT 468.930 245.720 469.930 247.850 ;
        RECT 470.770 245.720 471.770 247.850 ;
        RECT 472.610 245.720 473.610 247.850 ;
        RECT 474.450 245.720 475.450 247.850 ;
        RECT 476.290 245.720 477.290 247.850 ;
        RECT 478.130 245.720 479.130 247.850 ;
        RECT 479.970 245.720 480.970 247.850 ;
        RECT 481.810 245.720 482.810 247.850 ;
        RECT 483.650 245.720 484.650 247.850 ;
        RECT 485.490 245.720 486.490 247.850 ;
        RECT 487.330 245.720 488.330 247.850 ;
        RECT 489.170 245.720 490.170 247.850 ;
        RECT 491.010 245.720 492.010 247.850 ;
        RECT 492.850 245.720 493.850 247.850 ;
        RECT 494.690 245.720 495.690 247.850 ;
        RECT 496.530 245.720 497.530 247.850 ;
        RECT 498.370 245.720 499.370 247.850 ;
        RECT 500.210 245.720 501.210 247.850 ;
        RECT 502.050 245.720 503.050 247.850 ;
        RECT 503.890 245.720 504.890 247.850 ;
        RECT 505.730 245.720 506.730 247.850 ;
        RECT 507.570 245.720 508.570 247.850 ;
        RECT 509.410 245.720 510.410 247.850 ;
        RECT 511.250 245.720 512.250 247.850 ;
        RECT 513.090 245.720 514.090 247.850 ;
        RECT 514.930 245.720 515.930 247.850 ;
        RECT 516.770 245.720 517.770 247.850 ;
        RECT 518.610 245.720 519.610 247.850 ;
        RECT 520.450 245.720 521.450 247.850 ;
        RECT 522.290 245.720 523.290 247.850 ;
        RECT 524.130 245.720 525.130 247.850 ;
        RECT 525.970 245.720 526.970 247.850 ;
        RECT 527.810 245.720 528.810 247.850 ;
        RECT 529.650 245.720 530.650 247.850 ;
        RECT 531.490 245.720 532.490 247.850 ;
        RECT 533.330 245.720 534.330 247.850 ;
        RECT 535.170 245.720 536.170 247.850 ;
        RECT 537.010 245.720 538.010 247.850 ;
        RECT 538.850 245.720 539.850 247.850 ;
        RECT 540.690 245.720 541.690 247.850 ;
        RECT 542.530 245.720 543.530 247.850 ;
        RECT 544.370 245.720 545.370 247.850 ;
        RECT 546.210 245.720 547.210 247.850 ;
        RECT 548.050 245.720 549.050 247.850 ;
        RECT 549.890 245.720 550.890 247.850 ;
        RECT 551.730 245.720 552.730 247.850 ;
        RECT 553.570 245.720 554.570 247.850 ;
        RECT 555.410 245.720 556.410 247.850 ;
        RECT 557.250 245.720 558.250 247.850 ;
        RECT 559.090 245.720 560.090 247.850 ;
        RECT 560.930 245.720 561.930 247.850 ;
        RECT 562.770 245.720 563.770 247.850 ;
        RECT 564.610 245.720 565.610 247.850 ;
        RECT 566.450 245.720 567.450 247.850 ;
        RECT 568.290 245.720 569.290 247.850 ;
        RECT 570.130 245.720 571.130 247.850 ;
        RECT 571.970 245.720 572.970 247.850 ;
        RECT 573.810 245.720 574.810 247.850 ;
        RECT 575.650 245.720 576.650 247.850 ;
        RECT 577.490 245.720 578.490 247.850 ;
        RECT 579.330 245.720 580.330 247.850 ;
        RECT 581.170 245.720 582.170 247.850 ;
        RECT 583.010 245.720 584.010 247.850 ;
        RECT 584.850 245.720 585.850 247.850 ;
        RECT 586.690 245.720 587.690 247.850 ;
        RECT 588.530 245.720 589.530 247.850 ;
        RECT 590.370 245.720 591.370 247.850 ;
        RECT 592.210 245.720 593.210 247.850 ;
        RECT 594.050 245.720 595.050 247.850 ;
        RECT 595.890 245.720 596.890 247.850 ;
        RECT 597.730 245.720 598.730 247.850 ;
        RECT 599.570 245.720 600.570 247.850 ;
        RECT 601.410 245.720 602.410 247.850 ;
        RECT 603.250 245.720 643.440 247.850 ;
        RECT 0.100 4.280 643.440 245.720 ;
        RECT 0.100 0.010 26.490 4.280 ;
        RECT 27.330 0.010 32.010 4.280 ;
        RECT 32.850 0.010 37.530 4.280 ;
        RECT 38.370 0.010 43.050 4.280 ;
        RECT 43.890 0.010 48.570 4.280 ;
        RECT 49.410 0.010 54.090 4.280 ;
        RECT 54.930 0.010 59.610 4.280 ;
        RECT 60.450 0.010 65.130 4.280 ;
        RECT 65.970 0.010 70.650 4.280 ;
        RECT 71.490 0.010 76.170 4.280 ;
        RECT 77.010 0.010 81.690 4.280 ;
        RECT 82.530 0.010 87.210 4.280 ;
        RECT 88.050 0.010 92.730 4.280 ;
        RECT 93.570 0.010 98.250 4.280 ;
        RECT 99.090 0.010 103.770 4.280 ;
        RECT 104.610 0.010 109.290 4.280 ;
        RECT 110.130 0.010 114.810 4.280 ;
        RECT 115.650 0.010 120.330 4.280 ;
        RECT 121.170 0.010 125.850 4.280 ;
        RECT 126.690 0.010 131.370 4.280 ;
        RECT 132.210 0.010 136.890 4.280 ;
        RECT 137.730 0.010 142.410 4.280 ;
        RECT 143.250 0.010 147.930 4.280 ;
        RECT 148.770 0.010 153.450 4.280 ;
        RECT 154.290 0.010 158.970 4.280 ;
        RECT 159.810 0.010 164.490 4.280 ;
        RECT 165.330 0.010 170.010 4.280 ;
        RECT 170.850 0.010 175.530 4.280 ;
        RECT 176.370 0.010 181.050 4.280 ;
        RECT 181.890 0.010 186.570 4.280 ;
        RECT 187.410 0.010 192.090 4.280 ;
        RECT 192.930 0.010 197.610 4.280 ;
        RECT 198.450 0.010 203.130 4.280 ;
        RECT 203.970 0.010 208.650 4.280 ;
        RECT 209.490 0.010 214.170 4.280 ;
        RECT 215.010 0.010 219.690 4.280 ;
        RECT 220.530 0.010 225.210 4.280 ;
        RECT 226.050 0.010 230.730 4.280 ;
        RECT 231.570 0.010 236.250 4.280 ;
        RECT 237.090 0.010 241.770 4.280 ;
        RECT 242.610 0.010 247.290 4.280 ;
        RECT 248.130 0.010 252.810 4.280 ;
        RECT 253.650 0.010 258.330 4.280 ;
        RECT 259.170 0.010 263.850 4.280 ;
        RECT 264.690 0.010 269.370 4.280 ;
        RECT 270.210 0.010 274.890 4.280 ;
        RECT 275.730 0.010 280.410 4.280 ;
        RECT 281.250 0.010 285.930 4.280 ;
        RECT 286.770 0.010 291.450 4.280 ;
        RECT 292.290 0.010 296.970 4.280 ;
        RECT 297.810 0.010 302.490 4.280 ;
        RECT 303.330 0.010 308.010 4.280 ;
        RECT 308.850 0.010 313.530 4.280 ;
        RECT 314.370 0.010 319.050 4.280 ;
        RECT 319.890 0.010 324.570 4.280 ;
        RECT 325.410 0.010 330.090 4.280 ;
        RECT 330.930 0.010 335.610 4.280 ;
        RECT 336.450 0.010 341.130 4.280 ;
        RECT 341.970 0.010 346.650 4.280 ;
        RECT 347.490 0.010 352.170 4.280 ;
        RECT 353.010 0.010 357.690 4.280 ;
        RECT 358.530 0.010 363.210 4.280 ;
        RECT 364.050 0.010 368.730 4.280 ;
        RECT 369.570 0.010 374.250 4.280 ;
        RECT 375.090 0.010 379.770 4.280 ;
        RECT 380.610 0.010 385.290 4.280 ;
        RECT 386.130 0.010 390.810 4.280 ;
        RECT 391.650 0.010 396.330 4.280 ;
        RECT 397.170 0.010 401.850 4.280 ;
        RECT 402.690 0.010 407.370 4.280 ;
        RECT 408.210 0.010 412.890 4.280 ;
        RECT 413.730 0.010 418.410 4.280 ;
        RECT 419.250 0.010 423.930 4.280 ;
        RECT 424.770 0.010 429.450 4.280 ;
        RECT 430.290 0.010 434.970 4.280 ;
        RECT 435.810 0.010 440.490 4.280 ;
        RECT 441.330 0.010 446.010 4.280 ;
        RECT 446.850 0.010 451.530 4.280 ;
        RECT 452.370 0.010 457.050 4.280 ;
        RECT 457.890 0.010 462.570 4.280 ;
        RECT 463.410 0.010 468.090 4.280 ;
        RECT 468.930 0.010 473.610 4.280 ;
        RECT 474.450 0.010 479.130 4.280 ;
        RECT 479.970 0.010 484.650 4.280 ;
        RECT 485.490 0.010 490.170 4.280 ;
        RECT 491.010 0.010 495.690 4.280 ;
        RECT 496.530 0.010 501.210 4.280 ;
        RECT 502.050 0.010 506.730 4.280 ;
        RECT 507.570 0.010 512.250 4.280 ;
        RECT 513.090 0.010 517.770 4.280 ;
        RECT 518.610 0.010 523.290 4.280 ;
        RECT 524.130 0.010 528.810 4.280 ;
        RECT 529.650 0.010 534.330 4.280 ;
        RECT 535.170 0.010 539.850 4.280 ;
        RECT 540.690 0.010 545.370 4.280 ;
        RECT 546.210 0.010 550.890 4.280 ;
        RECT 551.730 0.010 556.410 4.280 ;
        RECT 557.250 0.010 561.930 4.280 ;
        RECT 562.770 0.010 567.450 4.280 ;
        RECT 568.290 0.010 572.970 4.280 ;
        RECT 573.810 0.010 578.490 4.280 ;
        RECT 579.330 0.010 584.010 4.280 ;
        RECT 584.850 0.010 589.530 4.280 ;
        RECT 590.370 0.010 595.050 4.280 ;
        RECT 595.890 0.010 600.570 4.280 ;
        RECT 601.410 0.010 606.090 4.280 ;
        RECT 606.930 0.010 611.610 4.280 ;
        RECT 612.450 0.010 617.130 4.280 ;
        RECT 617.970 0.010 622.650 4.280 ;
        RECT 623.490 0.010 643.440 4.280 ;
      LAYER met3 ;
        RECT 0.985 0.175 643.015 245.985 ;
      LAYER met4 ;
        RECT 1.215 237.280 640.945 245.305 ;
        RECT 1.215 182.880 20.640 237.280 ;
        RECT 1.215 10.240 7.540 182.880 ;
        RECT 9.940 10.240 10.300 182.880 ;
        RECT 12.700 178.760 20.640 182.880 ;
        RECT 23.040 178.760 97.440 237.280 ;
        RECT 99.840 178.760 174.240 237.280 ;
        RECT 176.640 178.760 251.040 237.280 ;
        RECT 253.440 178.760 327.840 237.280 ;
        RECT 330.240 178.760 404.640 237.280 ;
        RECT 407.040 178.760 481.440 237.280 ;
        RECT 483.840 178.760 558.240 237.280 ;
        RECT 560.640 180.160 635.040 237.280 ;
        RECT 560.640 178.760 630.380 180.160 ;
        RECT 12.700 10.240 630.380 178.760 ;
        RECT 632.780 10.240 635.040 180.160 ;
        RECT 637.440 10.240 640.945 237.280 ;
        RECT 1.215 0.175 640.945 10.240 ;
  END
END DataCache
END LIBRARY

