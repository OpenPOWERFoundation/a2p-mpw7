module SEL_PRI_32x4 (
  input      [31:0]   src0,
  input      [31:0]   src1,
  input      [31:0]   src2,
  input      [31:0]   src3,
  input      [3:0]    sel,
  output reg [31:0]   result
);
endmodule